magic
tech sky130A
magscale 1 2
timestamp 1665685787
<< error_p >>
rect -319 561 -295 673
rect -319 537 -154 561
rect -178 336 -154 537
<< rlocali >>
rect -353 537 -319 673
rect -353 503 -178 537
rect -212 336 -178 503
<< metal1 >>
rect 882 622 1192 698
rect 882 544 1012 622
rect 1100 544 1192 622
rect 882 442 1192 544
<< metal4 >>
rect 16 590 114 700
<< labels >>
flabel space 70 912 70 912 0 FreeSans 320 0 0 0 Exercise_3a
flabel space 64 828 64 828 0 FreeSans 320 0 0 0 Minimum_area_rule
flabel space 1042 944 1042 944 0 FreeSans 320 0 0 0 Exercise_3b
flabel space 1018 844 1018 844 0 FreeSans 320 0 0 0 Minimum_hole_rule
flabel space 1000 334 1000 334 0 FreeSans 320 0 0 0 *must_use_drc_style_sky130(full)*
<< end >>
