* NGSPICE file created from mgmt_protect.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
X0 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X2 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_193_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_193_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X19 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 VGND TE a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X24 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X28 Z A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X33 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt mprj2_logic_high HI vccd2 vssd2
XFILLER_0_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_170 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_71 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XPHY_0 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_1 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_30 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_2 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_207 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_1_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_112 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_59 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_170 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_129 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_199 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_187 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_100 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_112 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_146 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_158 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_71 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
Xinst vssd2 vssd2 vccd2 vccd2 HI inst/LO sky130_fd_sc_hd__conb_1
XFILLER_0_117 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_129 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_30 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_42 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_204 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_8
XFILLER_0_54 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_88 vssd2 vssd2 vccd2 vccd2 sky130_fd_sc_hd__decap_12
.ends

.subckt mprj_logic_high HI[199] HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105]
+ HI[106] HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115]
+ HI[116] HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125]
+ HI[126] HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135]
+ HI[136] HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145]
+ HI[146] HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155]
+ HI[156] HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165]
+ HI[166] HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175]
+ HI[176] HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185]
+ HI[186] HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195]
+ HI[196] HI[197] HI[198] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[46] HI[47]
+ HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57] HI[58]
+ HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68] HI[69]
+ HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79] HI[7]
+ HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8] HI[90]
+ HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1 vssd1
+
Xinsts\[308\] vssd1 vssd1 vccd1 vccd1 HI[308] insts\[308\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[210\] vssd1 vssd1 vccd1 vccd1 HI[210] insts\[210\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[425\] vssd1 vssd1 vccd1 vccd1 HI[425] insts\[425\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[258\] vssd1 vssd1 vccd1 vccd1 HI[258] insts\[258\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[160\] vssd1 vssd1 vccd1 vccd1 HI[160] insts\[160\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[40\] vssd1 vssd1 vccd1 vccd1 HI[40] insts\[40\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[375\] vssd1 vssd1 vccd1 vccd1 HI[375] insts\[375\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[88\] vssd1 vssd1 vccd1 vccd1 HI[88] insts\[88\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[123\] vssd1 vssd1 vccd1 vccd1 HI[123] insts\[123\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[240\] vssd1 vssd1 vccd1 vccd1 HI[240] insts\[240\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[338\] vssd1 vssd1 vccd1 vccd1 HI[338] insts\[338\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[9\] vssd1 vssd1 vccd1 vccd1 HI[9] insts\[9\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[455\] vssd1 vssd1 vccd1 vccd1 HI[455] insts\[455\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[288\] vssd1 vssd1 vccd1 vccd1 HI[288] insts\[288\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[190\] vssd1 vssd1 vccd1 vccd1 HI[190] insts\[190\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[70\] vssd1 vssd1 vccd1 vccd1 HI[70] insts\[70\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[203\] vssd1 vssd1 vccd1 vccd1 HI[203] insts\[203\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[418\] vssd1 vssd1 vccd1 vccd1 HI[418] insts\[418\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[153\] vssd1 vssd1 vccd1 vccd1 HI[153] insts\[153\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[320\] vssd1 vssd1 vccd1 vccd1 HI[320] insts\[320\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[33\] vssd1 vssd1 vccd1 vccd1 HI[33] insts\[33\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[270\] vssd1 vssd1 vccd1 vccd1 HI[270] insts\[270\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[368\] vssd1 vssd1 vccd1 vccd1 HI[368] insts\[368\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[116\] vssd1 vssd1 vccd1 vccd1 HI[116] insts\[116\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[233\] vssd1 vssd1 vccd1 vccd1 HI[233] insts\[233\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[400\] vssd1 vssd1 vccd1 vccd1 HI[400] insts\[400\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[183\] vssd1 vssd1 vccd1 vccd1 HI[183] insts\[183\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[448\] vssd1 vssd1 vccd1 vccd1 HI[448] insts\[448\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[350\] vssd1 vssd1 vccd1 vccd1 HI[350] insts\[350\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[63\] vssd1 vssd1 vccd1 vccd1 HI[63] insts\[63\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[398\] vssd1 vssd1 vccd1 vccd1 HI[398] insts\[398\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[146\] vssd1 vssd1 vccd1 vccd1 HI[146] insts\[146\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[313\] vssd1 vssd1 vccd1 vccd1 HI[313] insts\[313\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[26\] vssd1 vssd1 vccd1 vccd1 HI[26] insts\[26\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[430\] vssd1 vssd1 vccd1 vccd1 HI[430] insts\[430\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[263\] vssd1 vssd1 vccd1 vccd1 HI[263] insts\[263\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[109\] vssd1 vssd1 vccd1 vccd1 HI[109] insts\[109\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[380\] vssd1 vssd1 vccd1 vccd1 HI[380] insts\[380\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[93\] vssd1 vssd1 vccd1 vccd1 HI[93] insts\[93\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[226\] vssd1 vssd1 vccd1 vccd1 HI[226] insts\[226\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[343\] vssd1 vssd1 vccd1 vccd1 HI[343] insts\[343\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[176\] vssd1 vssd1 vccd1 vccd1 HI[176] insts\[176\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[56\] vssd1 vssd1 vccd1 vccd1 HI[56] insts\[56\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[460\] vssd1 vssd1 vccd1 vccd1 HI[460] insts\[460\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[293\] vssd1 vssd1 vccd1 vccd1 HI[293] insts\[293\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[139\] vssd1 vssd1 vccd1 vccd1 HI[139] insts\[139\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[306\] vssd1 vssd1 vccd1 vccd1 HI[306] insts\[306\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[19\] vssd1 vssd1 vccd1 vccd1 HI[19] insts\[19\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[423\] vssd1 vssd1 vccd1 vccd1 HI[423] insts\[423\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[256\] vssd1 vssd1 vccd1 vccd1 HI[256] insts\[256\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[373\] vssd1 vssd1 vccd1 vccd1 HI[373] insts\[373\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[86\] vssd1 vssd1 vccd1 vccd1 HI[86] insts\[86\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[219\] vssd1 vssd1 vccd1 vccd1 HI[219] insts\[219\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[121\] vssd1 vssd1 vccd1 vccd1 HI[121] insts\[121\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[336\] vssd1 vssd1 vccd1 vccd1 HI[336] insts\[336\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[169\] vssd1 vssd1 vccd1 vccd1 HI[169] insts\[169\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[49\] vssd1 vssd1 vccd1 vccd1 HI[49] insts\[49\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[286\] vssd1 vssd1 vccd1 vccd1 HI[286] insts\[286\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[7\] vssd1 vssd1 vccd1 vccd1 HI[7] insts\[7\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[453\] vssd1 vssd1 vccd1 vccd1 HI[453] insts\[453\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[201\] vssd1 vssd1 vccd1 vccd1 HI[201] insts\[201\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[416\] vssd1 vssd1 vccd1 vccd1 HI[416] insts\[416\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[249\] vssd1 vssd1 vccd1 vccd1 HI[249] insts\[249\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[151\] vssd1 vssd1 vccd1 vccd1 HI[151] insts\[151\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[31\] vssd1 vssd1 vccd1 vccd1 HI[31] insts\[31\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[199\] vssd1 vssd1 vccd1 vccd1 HI[199] insts\[199\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[366\] vssd1 vssd1 vccd1 vccd1 HI[366] insts\[366\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[79\] vssd1 vssd1 vccd1 vccd1 HI[79] insts\[79\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[114\] vssd1 vssd1 vccd1 vccd1 HI[114] insts\[114\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[231\] vssd1 vssd1 vccd1 vccd1 HI[231] insts\[231\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[329\] vssd1 vssd1 vccd1 vccd1 HI[329] insts\[329\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[446\] vssd1 vssd1 vccd1 vccd1 HI[446] insts\[446\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[279\] vssd1 vssd1 vccd1 vccd1 HI[279] insts\[279\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[181\] vssd1 vssd1 vccd1 vccd1 HI[181] insts\[181\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[61\] vssd1 vssd1 vccd1 vccd1 HI[61] insts\[61\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[396\] vssd1 vssd1 vccd1 vccd1 HI[396] insts\[396\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[144\] vssd1 vssd1 vccd1 vccd1 HI[144] insts\[144\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[311\] vssd1 vssd1 vccd1 vccd1 HI[311] insts\[311\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[409\] vssd1 vssd1 vccd1 vccd1 HI[409] insts\[409\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[24\] vssd1 vssd1 vccd1 vccd1 HI[24] insts\[24\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[261\] vssd1 vssd1 vccd1 vccd1 HI[261] insts\[261\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[359\] vssd1 vssd1 vccd1 vccd1 HI[359] insts\[359\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[107\] vssd1 vssd1 vccd1 vccd1 HI[107] insts\[107\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[91\] vssd1 vssd1 vccd1 vccd1 HI[91] insts\[91\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[224\] vssd1 vssd1 vccd1 vccd1 HI[224] insts\[224\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[439\] vssd1 vssd1 vccd1 vccd1 HI[439] insts\[439\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[174\] vssd1 vssd1 vccd1 vccd1 HI[174] insts\[174\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[341\] vssd1 vssd1 vccd1 vccd1 HI[341] insts\[341\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[54\] vssd1 vssd1 vccd1 vccd1 HI[54] insts\[54\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[291\] vssd1 vssd1 vccd1 vccd1 HI[291] insts\[291\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[389\] vssd1 vssd1 vccd1 vccd1 HI[389] insts\[389\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[304\] vssd1 vssd1 vccd1 vccd1 HI[304] insts\[304\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[137\] vssd1 vssd1 vccd1 vccd1 HI[137] insts\[137\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[17\] vssd1 vssd1 vccd1 vccd1 HI[17] insts\[17\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[421\] vssd1 vssd1 vccd1 vccd1 HI[421] insts\[421\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[254\] vssd1 vssd1 vccd1 vccd1 HI[254] insts\[254\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[371\] vssd1 vssd1 vccd1 vccd1 HI[371] insts\[371\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[84\] vssd1 vssd1 vccd1 vccd1 HI[84] insts\[84\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[217\] vssd1 vssd1 vccd1 vccd1 HI[217] insts\[217\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[167\] vssd1 vssd1 vccd1 vccd1 HI[167] insts\[167\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[334\] vssd1 vssd1 vccd1 vccd1 HI[334] insts\[334\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[47\] vssd1 vssd1 vccd1 vccd1 HI[47] insts\[47\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[5\] vssd1 vssd1 vccd1 vccd1 HI[5] insts\[5\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[451\] vssd1 vssd1 vccd1 vccd1 HI[451] insts\[451\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[284\] vssd1 vssd1 vccd1 vccd1 HI[284] insts\[284\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[247\] vssd1 vssd1 vccd1 vccd1 HI[247] insts\[247\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[414\] vssd1 vssd1 vccd1 vccd1 HI[414] insts\[414\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[197\] vssd1 vssd1 vccd1 vccd1 HI[197] insts\[197\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[364\] vssd1 vssd1 vccd1 vccd1 HI[364] insts\[364\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[77\] vssd1 vssd1 vccd1 vccd1 HI[77] insts\[77\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[112\] vssd1 vssd1 vccd1 vccd1 HI[112] insts\[112\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[327\] vssd1 vssd1 vccd1 vccd1 HI[327] insts\[327\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[444\] vssd1 vssd1 vccd1 vccd1 HI[444] insts\[444\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[277\] vssd1 vssd1 vccd1 vccd1 HI[277] insts\[277\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[394\] vssd1 vssd1 vccd1 vccd1 HI[394] insts\[394\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[407\] vssd1 vssd1 vccd1 vccd1 HI[407] insts\[407\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[142\] vssd1 vssd1 vccd1 vccd1 HI[142] insts\[142\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[22\] vssd1 vssd1 vccd1 vccd1 HI[22] insts\[22\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[357\] vssd1 vssd1 vccd1 vccd1 HI[357] insts\[357\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[105\] vssd1 vssd1 vccd1 vccd1 HI[105] insts\[105\]/LO sky130_fd_sc_hd__conb_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[222\] vssd1 vssd1 vccd1 vccd1 HI[222] insts\[222\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[437\] vssd1 vssd1 vccd1 vccd1 HI[437] insts\[437\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[172\] vssd1 vssd1 vccd1 vccd1 HI[172] insts\[172\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[52\] vssd1 vssd1 vccd1 vccd1 HI[52] insts\[52\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[387\] vssd1 vssd1 vccd1 vccd1 HI[387] insts\[387\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[302\] vssd1 vssd1 vccd1 vccd1 HI[302] insts\[302\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[135\] vssd1 vssd1 vccd1 vccd1 HI[135] insts\[135\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[15\] vssd1 vssd1 vccd1 vccd1 HI[15] insts\[15\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[252\] vssd1 vssd1 vccd1 vccd1 HI[252] insts\[252\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[82\] vssd1 vssd1 vccd1 vccd1 HI[82] insts\[82\]/LO sky130_fd_sc_hd__conb_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[215\] vssd1 vssd1 vccd1 vccd1 HI[215] insts\[215\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[165\] vssd1 vssd1 vccd1 vccd1 HI[165] insts\[165\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[332\] vssd1 vssd1 vccd1 vccd1 HI[332] insts\[332\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[45\] vssd1 vssd1 vccd1 vccd1 HI[45] insts\[45\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[282\] vssd1 vssd1 vccd1 vccd1 HI[282] insts\[282\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[3\] vssd1 vssd1 vccd1 vccd1 HI[3] insts\[3\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[128\] vssd1 vssd1 vccd1 vccd1 HI[128] insts\[128\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[245\] vssd1 vssd1 vccd1 vccd1 HI[245] insts\[245\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[412\] vssd1 vssd1 vccd1 vccd1 HI[412] insts\[412\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[195\] vssd1 vssd1 vccd1 vccd1 HI[195] insts\[195\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[362\] vssd1 vssd1 vccd1 vccd1 HI[362] insts\[362\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[75\] vssd1 vssd1 vccd1 vccd1 HI[75] insts\[75\]/LO sky130_fd_sc_hd__conb_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[208\] vssd1 vssd1 vccd1 vccd1 HI[208] insts\[208\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[110\] vssd1 vssd1 vccd1 vccd1 HI[110] insts\[110\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[158\] vssd1 vssd1 vccd1 vccd1 HI[158] insts\[158\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[325\] vssd1 vssd1 vccd1 vccd1 HI[325] insts\[325\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[38\] vssd1 vssd1 vccd1 vccd1 HI[38] insts\[38\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[442\] vssd1 vssd1 vccd1 vccd1 HI[442] insts\[442\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[275\] vssd1 vssd1 vccd1 vccd1 HI[275] insts\[275\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[392\] vssd1 vssd1 vccd1 vccd1 HI[392] insts\[392\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[238\] vssd1 vssd1 vccd1 vccd1 HI[238] insts\[238\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[140\] vssd1 vssd1 vccd1 vccd1 HI[140] insts\[140\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[405\] vssd1 vssd1 vccd1 vccd1 HI[405] insts\[405\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[20\] vssd1 vssd1 vccd1 vccd1 HI[20] insts\[20\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[188\] vssd1 vssd1 vccd1 vccd1 HI[188] insts\[188\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[355\] vssd1 vssd1 vccd1 vccd1 HI[355] insts\[355\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[68\] vssd1 vssd1 vccd1 vccd1 HI[68] insts\[68\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[103\] vssd1 vssd1 vccd1 vccd1 HI[103] insts\[103\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[220\] vssd1 vssd1 vccd1 vccd1 HI[220] insts\[220\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[318\] vssd1 vssd1 vccd1 vccd1 HI[318] insts\[318\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[170\] vssd1 vssd1 vccd1 vccd1 HI[170] insts\[170\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[435\] vssd1 vssd1 vccd1 vccd1 HI[435] insts\[435\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[268\] vssd1 vssd1 vccd1 vccd1 HI[268] insts\[268\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[50\] vssd1 vssd1 vccd1 vccd1 HI[50] insts\[50\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[385\] vssd1 vssd1 vccd1 vccd1 HI[385] insts\[385\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[98\] vssd1 vssd1 vccd1 vccd1 HI[98] insts\[98\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[300\] vssd1 vssd1 vccd1 vccd1 HI[300] insts\[300\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[133\] vssd1 vssd1 vccd1 vccd1 HI[133] insts\[133\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[13\] vssd1 vssd1 vccd1 vccd1 HI[13] insts\[13\]/LO sky130_fd_sc_hd__conb_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[250\] vssd1 vssd1 vccd1 vccd1 HI[250] insts\[250\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[348\] vssd1 vssd1 vccd1 vccd1 HI[348] insts\[348\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[298\] vssd1 vssd1 vccd1 vccd1 HI[298] insts\[298\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[80\] vssd1 vssd1 vccd1 vccd1 HI[80] insts\[80\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[213\] vssd1 vssd1 vccd1 vccd1 HI[213] insts\[213\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[428\] vssd1 vssd1 vccd1 vccd1 HI[428] insts\[428\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[163\] vssd1 vssd1 vccd1 vccd1 HI[163] insts\[163\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[330\] vssd1 vssd1 vccd1 vccd1 HI[330] insts\[330\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[43\] vssd1 vssd1 vccd1 vccd1 HI[43] insts\[43\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[280\] vssd1 vssd1 vccd1 vccd1 HI[280] insts\[280\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[1\] vssd1 vssd1 vccd1 vccd1 HI[1] insts\[1\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[378\] vssd1 vssd1 vccd1 vccd1 HI[378] insts\[378\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[126\] vssd1 vssd1 vccd1 vccd1 HI[126] insts\[126\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[243\] vssd1 vssd1 vccd1 vccd1 HI[243] insts\[243\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[410\] vssd1 vssd1 vccd1 vccd1 HI[410] insts\[410\]/LO sky130_fd_sc_hd__conb_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[458\] vssd1 vssd1 vccd1 vccd1 HI[458] insts\[458\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[193\] vssd1 vssd1 vccd1 vccd1 HI[193] insts\[193\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[360\] vssd1 vssd1 vccd1 vccd1 HI[360] insts\[360\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[73\] vssd1 vssd1 vccd1 vccd1 HI[73] insts\[73\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[206\] vssd1 vssd1 vccd1 vccd1 HI[206] insts\[206\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[156\] vssd1 vssd1 vccd1 vccd1 HI[156] insts\[156\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[323\] vssd1 vssd1 vccd1 vccd1 HI[323] insts\[323\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[36\] vssd1 vssd1 vccd1 vccd1 HI[36] insts\[36\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[273\] vssd1 vssd1 vccd1 vccd1 HI[273] insts\[273\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[440\] vssd1 vssd1 vccd1 vccd1 HI[440] insts\[440\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[119\] vssd1 vssd1 vccd1 vccd1 HI[119] insts\[119\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[390\] vssd1 vssd1 vccd1 vccd1 HI[390] insts\[390\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[236\] vssd1 vssd1 vccd1 vccd1 HI[236] insts\[236\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[403\] vssd1 vssd1 vccd1 vccd1 HI[403] insts\[403\]/LO sky130_fd_sc_hd__conb_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[353\] vssd1 vssd1 vccd1 vccd1 HI[353] insts\[353\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[186\] vssd1 vssd1 vccd1 vccd1 HI[186] insts\[186\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[66\] vssd1 vssd1 vccd1 vccd1 HI[66] insts\[66\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[101\] vssd1 vssd1 vccd1 vccd1 HI[101] insts\[101\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[316\] vssd1 vssd1 vccd1 vccd1 HI[316] insts\[316\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[149\] vssd1 vssd1 vccd1 vccd1 HI[149] insts\[149\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[29\] vssd1 vssd1 vccd1 vccd1 HI[29] insts\[29\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[433\] vssd1 vssd1 vccd1 vccd1 HI[433] insts\[433\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[266\] vssd1 vssd1 vccd1 vccd1 HI[266] insts\[266\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[383\] vssd1 vssd1 vccd1 vccd1 HI[383] insts\[383\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[96\] vssd1 vssd1 vccd1 vccd1 HI[96] insts\[96\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[229\] vssd1 vssd1 vccd1 vccd1 HI[229] insts\[229\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[131\] vssd1 vssd1 vccd1 vccd1 HI[131] insts\[131\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[11\] vssd1 vssd1 vccd1 vccd1 HI[11] insts\[11\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[179\] vssd1 vssd1 vccd1 vccd1 HI[179] insts\[179\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[346\] vssd1 vssd1 vccd1 vccd1 HI[346] insts\[346\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[59\] vssd1 vssd1 vccd1 vccd1 HI[59] insts\[59\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[296\] vssd1 vssd1 vccd1 vccd1 HI[296] insts\[296\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[211\] vssd1 vssd1 vccd1 vccd1 HI[211] insts\[211\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[309\] vssd1 vssd1 vccd1 vccd1 HI[309] insts\[309\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[426\] vssd1 vssd1 vccd1 vccd1 HI[426] insts\[426\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[259\] vssd1 vssd1 vccd1 vccd1 HI[259] insts\[259\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[161\] vssd1 vssd1 vccd1 vccd1 HI[161] insts\[161\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[41\] vssd1 vssd1 vccd1 vccd1 HI[41] insts\[41\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[376\] vssd1 vssd1 vccd1 vccd1 HI[376] insts\[376\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[89\] vssd1 vssd1 vccd1 vccd1 HI[89] insts\[89\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[124\] vssd1 vssd1 vccd1 vccd1 HI[124] insts\[124\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[241\] vssd1 vssd1 vccd1 vccd1 HI[241] insts\[241\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[339\] vssd1 vssd1 vccd1 vccd1 HI[339] insts\[339\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[456\] vssd1 vssd1 vccd1 vccd1 HI[456] insts\[456\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[289\] vssd1 vssd1 vccd1 vccd1 HI[289] insts\[289\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[191\] vssd1 vssd1 vccd1 vccd1 HI[191] insts\[191\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[71\] vssd1 vssd1 vccd1 vccd1 HI[71] insts\[71\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[204\] vssd1 vssd1 vccd1 vccd1 HI[204] insts\[204\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[419\] vssd1 vssd1 vccd1 vccd1 HI[419] insts\[419\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[154\] vssd1 vssd1 vccd1 vccd1 HI[154] insts\[154\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[321\] vssd1 vssd1 vccd1 vccd1 HI[321] insts\[321\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[34\] vssd1 vssd1 vccd1 vccd1 HI[34] insts\[34\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[271\] vssd1 vssd1 vccd1 vccd1 HI[271] insts\[271\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[369\] vssd1 vssd1 vccd1 vccd1 HI[369] insts\[369\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[117\] vssd1 vssd1 vccd1 vccd1 HI[117] insts\[117\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[234\] vssd1 vssd1 vccd1 vccd1 HI[234] insts\[234\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[401\] vssd1 vssd1 vccd1 vccd1 HI[401] insts\[401\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[449\] vssd1 vssd1 vccd1 vccd1 HI[449] insts\[449\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[184\] vssd1 vssd1 vccd1 vccd1 HI[184] insts\[184\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[351\] vssd1 vssd1 vccd1 vccd1 HI[351] insts\[351\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[64\] vssd1 vssd1 vccd1 vccd1 HI[64] insts\[64\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[399\] vssd1 vssd1 vccd1 vccd1 HI[399] insts\[399\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[314\] vssd1 vssd1 vccd1 vccd1 HI[314] insts\[314\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[147\] vssd1 vssd1 vccd1 vccd1 HI[147] insts\[147\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[27\] vssd1 vssd1 vccd1 vccd1 HI[27] insts\[27\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[431\] vssd1 vssd1 vccd1 vccd1 HI[431] insts\[431\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[264\] vssd1 vssd1 vccd1 vccd1 HI[264] insts\[264\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[381\] vssd1 vssd1 vccd1 vccd1 HI[381] insts\[381\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[94\] vssd1 vssd1 vccd1 vccd1 HI[94] insts\[94\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[227\] vssd1 vssd1 vccd1 vccd1 HI[227] insts\[227\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[177\] vssd1 vssd1 vccd1 vccd1 HI[177] insts\[177\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[344\] vssd1 vssd1 vccd1 vccd1 HI[344] insts\[344\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[57\] vssd1 vssd1 vccd1 vccd1 HI[57] insts\[57\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[461\] vssd1 vssd1 vccd1 vccd1 HI[461] insts\[461\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[294\] vssd1 vssd1 vccd1 vccd1 HI[294] insts\[294\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[307\] vssd1 vssd1 vccd1 vccd1 HI[307] insts\[307\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[424\] vssd1 vssd1 vccd1 vccd1 HI[424] insts\[424\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[257\] vssd1 vssd1 vccd1 vccd1 HI[257] insts\[257\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[374\] vssd1 vssd1 vccd1 vccd1 HI[374] insts\[374\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[87\] vssd1 vssd1 vccd1 vccd1 HI[87] insts\[87\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[122\] vssd1 vssd1 vccd1 vccd1 HI[122] insts\[122\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[337\] vssd1 vssd1 vccd1 vccd1 HI[337] insts\[337\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[8\] vssd1 vssd1 vccd1 vccd1 HI[8] insts\[8\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[454\] vssd1 vssd1 vccd1 vccd1 HI[454] insts\[454\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[287\] vssd1 vssd1 vccd1 vccd1 HI[287] insts\[287\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[202\] vssd1 vssd1 vccd1 vccd1 HI[202] insts\[202\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[417\] vssd1 vssd1 vccd1 vccd1 HI[417] insts\[417\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[152\] vssd1 vssd1 vccd1 vccd1 HI[152] insts\[152\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[32\] vssd1 vssd1 vccd1 vccd1 HI[32] insts\[32\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[367\] vssd1 vssd1 vccd1 vccd1 HI[367] insts\[367\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[115\] vssd1 vssd1 vccd1 vccd1 HI[115] insts\[115\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[232\] vssd1 vssd1 vccd1 vccd1 HI[232] insts\[232\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[447\] vssd1 vssd1 vccd1 vccd1 HI[447] insts\[447\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[182\] vssd1 vssd1 vccd1 vccd1 HI[182] insts\[182\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[62\] vssd1 vssd1 vccd1 vccd1 HI[62] insts\[62\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[397\] vssd1 vssd1 vccd1 vccd1 HI[397] insts\[397\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[145\] vssd1 vssd1 vccd1 vccd1 HI[145] insts\[145\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[312\] vssd1 vssd1 vccd1 vccd1 HI[312] insts\[312\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[25\] vssd1 vssd1 vccd1 vccd1 HI[25] insts\[25\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[262\] vssd1 vssd1 vccd1 vccd1 HI[262] insts\[262\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[108\] vssd1 vssd1 vccd1 vccd1 HI[108] insts\[108\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[92\] vssd1 vssd1 vccd1 vccd1 HI[92] insts\[92\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[225\] vssd1 vssd1 vccd1 vccd1 HI[225] insts\[225\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[175\] vssd1 vssd1 vccd1 vccd1 HI[175] insts\[175\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[342\] vssd1 vssd1 vccd1 vccd1 HI[342] insts\[342\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[55\] vssd1 vssd1 vccd1 vccd1 HI[55] insts\[55\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[292\] vssd1 vssd1 vccd1 vccd1 HI[292] insts\[292\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[305\] vssd1 vssd1 vccd1 vccd1 HI[305] insts\[305\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[138\] vssd1 vssd1 vccd1 vccd1 HI[138] insts\[138\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[18\] vssd1 vssd1 vccd1 vccd1 HI[18] insts\[18\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[422\] vssd1 vssd1 vccd1 vccd1 HI[422] insts\[422\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[255\] vssd1 vssd1 vccd1 vccd1 HI[255] insts\[255\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[372\] vssd1 vssd1 vccd1 vccd1 HI[372] insts\[372\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[85\] vssd1 vssd1 vccd1 vccd1 HI[85] insts\[85\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[218\] vssd1 vssd1 vccd1 vccd1 HI[218] insts\[218\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[120\] vssd1 vssd1 vccd1 vccd1 HI[120] insts\[120\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[168\] vssd1 vssd1 vccd1 vccd1 HI[168] insts\[168\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[335\] vssd1 vssd1 vccd1 vccd1 HI[335] insts\[335\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[48\] vssd1 vssd1 vccd1 vccd1 HI[48] insts\[48\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[6\] vssd1 vssd1 vccd1 vccd1 HI[6] insts\[6\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[452\] vssd1 vssd1 vccd1 vccd1 HI[452] insts\[452\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[285\] vssd1 vssd1 vccd1 vccd1 HI[285] insts\[285\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[200\] vssd1 vssd1 vccd1 vccd1 HI[200] insts\[200\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[415\] vssd1 vssd1 vccd1 vccd1 HI[415] insts\[415\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[248\] vssd1 vssd1 vccd1 vccd1 HI[248] insts\[248\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[150\] vssd1 vssd1 vccd1 vccd1 HI[150] insts\[150\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[30\] vssd1 vssd1 vccd1 vccd1 HI[30] insts\[30\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[198\] vssd1 vssd1 vccd1 vccd1 HI[198] insts\[198\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[365\] vssd1 vssd1 vccd1 vccd1 HI[365] insts\[365\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[78\] vssd1 vssd1 vccd1 vccd1 HI[78] insts\[78\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[113\] vssd1 vssd1 vccd1 vccd1 HI[113] insts\[113\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[230\] vssd1 vssd1 vccd1 vccd1 HI[230] insts\[230\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[328\] vssd1 vssd1 vccd1 vccd1 HI[328] insts\[328\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[445\] vssd1 vssd1 vccd1 vccd1 HI[445] insts\[445\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[278\] vssd1 vssd1 vccd1 vccd1 HI[278] insts\[278\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[180\] vssd1 vssd1 vccd1 vccd1 HI[180] insts\[180\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[60\] vssd1 vssd1 vccd1 vccd1 HI[60] insts\[60\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[395\] vssd1 vssd1 vccd1 vccd1 HI[395] insts\[395\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[310\] vssd1 vssd1 vccd1 vccd1 HI[310] insts\[310\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[143\] vssd1 vssd1 vccd1 vccd1 HI[143] insts\[143\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[408\] vssd1 vssd1 vccd1 vccd1 HI[408] insts\[408\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[23\] vssd1 vssd1 vccd1 vccd1 HI[23] insts\[23\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[260\] vssd1 vssd1 vccd1 vccd1 HI[260] insts\[260\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[358\] vssd1 vssd1 vccd1 vccd1 HI[358] insts\[358\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[106\] vssd1 vssd1 vccd1 vccd1 HI[106] insts\[106\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[90\] vssd1 vssd1 vccd1 vccd1 HI[90] insts\[90\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[223\] vssd1 vssd1 vccd1 vccd1 HI[223] insts\[223\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[438\] vssd1 vssd1 vccd1 vccd1 HI[438] insts\[438\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[173\] vssd1 vssd1 vccd1 vccd1 HI[173] insts\[173\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[340\] vssd1 vssd1 vccd1 vccd1 HI[340] insts\[340\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[53\] vssd1 vssd1 vccd1 vccd1 HI[53] insts\[53\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[290\] vssd1 vssd1 vccd1 vccd1 HI[290] insts\[290\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[388\] vssd1 vssd1 vccd1 vccd1 HI[388] insts\[388\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[303\] vssd1 vssd1 vccd1 vccd1 HI[303] insts\[303\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[136\] vssd1 vssd1 vccd1 vccd1 HI[136] insts\[136\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[16\] vssd1 vssd1 vccd1 vccd1 HI[16] insts\[16\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[420\] vssd1 vssd1 vccd1 vccd1 HI[420] insts\[420\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[253\] vssd1 vssd1 vccd1 vccd1 HI[253] insts\[253\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[370\] vssd1 vssd1 vccd1 vccd1 HI[370] insts\[370\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[83\] vssd1 vssd1 vccd1 vccd1 HI[83] insts\[83\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[216\] vssd1 vssd1 vccd1 vccd1 HI[216] insts\[216\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[166\] vssd1 vssd1 vccd1 vccd1 HI[166] insts\[166\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[333\] vssd1 vssd1 vccd1 vccd1 HI[333] insts\[333\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[46\] vssd1 vssd1 vccd1 vccd1 HI[46] insts\[46\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[450\] vssd1 vssd1 vccd1 vccd1 HI[450] insts\[450\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[283\] vssd1 vssd1 vccd1 vccd1 HI[283] insts\[283\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[4\] vssd1 vssd1 vccd1 vccd1 HI[4] insts\[4\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[129\] vssd1 vssd1 vccd1 vccd1 HI[129] insts\[129\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[413\] vssd1 vssd1 vccd1 vccd1 HI[413] insts\[413\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[246\] vssd1 vssd1 vccd1 vccd1 HI[246] insts\[246\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[196\] vssd1 vssd1 vccd1 vccd1 HI[196] insts\[196\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[363\] vssd1 vssd1 vccd1 vccd1 HI[363] insts\[363\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[76\] vssd1 vssd1 vccd1 vccd1 HI[76] insts\[76\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[209\] vssd1 vssd1 vccd1 vccd1 HI[209] insts\[209\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[111\] vssd1 vssd1 vccd1 vccd1 HI[111] insts\[111\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[159\] vssd1 vssd1 vccd1 vccd1 HI[159] insts\[159\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[326\] vssd1 vssd1 vccd1 vccd1 HI[326] insts\[326\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[39\] vssd1 vssd1 vccd1 vccd1 HI[39] insts\[39\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[443\] vssd1 vssd1 vccd1 vccd1 HI[443] insts\[443\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[276\] vssd1 vssd1 vccd1 vccd1 HI[276] insts\[276\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[393\] vssd1 vssd1 vccd1 vccd1 HI[393] insts\[393\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[239\] vssd1 vssd1 vccd1 vccd1 HI[239] insts\[239\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[141\] vssd1 vssd1 vccd1 vccd1 HI[141] insts\[141\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[406\] vssd1 vssd1 vccd1 vccd1 HI[406] insts\[406\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[21\] vssd1 vssd1 vccd1 vccd1 HI[21] insts\[21\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[189\] vssd1 vssd1 vccd1 vccd1 HI[189] insts\[189\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[356\] vssd1 vssd1 vccd1 vccd1 HI[356] insts\[356\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[69\] vssd1 vssd1 vccd1 vccd1 HI[69] insts\[69\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[104\] vssd1 vssd1 vccd1 vccd1 HI[104] insts\[104\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[221\] vssd1 vssd1 vccd1 vccd1 HI[221] insts\[221\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[319\] vssd1 vssd1 vccd1 vccd1 HI[319] insts\[319\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[436\] vssd1 vssd1 vccd1 vccd1 HI[436] insts\[436\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[269\] vssd1 vssd1 vccd1 vccd1 HI[269] insts\[269\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[171\] vssd1 vssd1 vccd1 vccd1 HI[171] insts\[171\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[51\] vssd1 vssd1 vccd1 vccd1 HI[51] insts\[51\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[386\] vssd1 vssd1 vccd1 vccd1 HI[386] insts\[386\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[99\] vssd1 vssd1 vccd1 vccd1 HI[99] insts\[99\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[301\] vssd1 vssd1 vccd1 vccd1 HI[301] insts\[301\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[134\] vssd1 vssd1 vccd1 vccd1 HI[134] insts\[134\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[14\] vssd1 vssd1 vccd1 vccd1 HI[14] insts\[14\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[251\] vssd1 vssd1 vccd1 vccd1 HI[251] insts\[251\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[349\] vssd1 vssd1 vccd1 vccd1 HI[349] insts\[349\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[299\] vssd1 vssd1 vccd1 vccd1 HI[299] insts\[299\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[81\] vssd1 vssd1 vccd1 vccd1 HI[81] insts\[81\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[214\] vssd1 vssd1 vccd1 vccd1 HI[214] insts\[214\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[429\] vssd1 vssd1 vccd1 vccd1 HI[429] insts\[429\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[164\] vssd1 vssd1 vccd1 vccd1 HI[164] insts\[164\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[331\] vssd1 vssd1 vccd1 vccd1 HI[331] insts\[331\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[44\] vssd1 vssd1 vccd1 vccd1 HI[44] insts\[44\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[2\] vssd1 vssd1 vccd1 vccd1 HI[2] insts\[2\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[281\] vssd1 vssd1 vccd1 vccd1 HI[281] insts\[281\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[379\] vssd1 vssd1 vccd1 vccd1 HI[379] insts\[379\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[127\] vssd1 vssd1 vccd1 vccd1 HI[127] insts\[127\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[244\] vssd1 vssd1 vccd1 vccd1 HI[244] insts\[244\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[411\] vssd1 vssd1 vccd1 vccd1 HI[411] insts\[411\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[459\] vssd1 vssd1 vccd1 vccd1 HI[459] insts\[459\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[194\] vssd1 vssd1 vccd1 vccd1 HI[194] insts\[194\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[361\] vssd1 vssd1 vccd1 vccd1 HI[361] insts\[361\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[74\] vssd1 vssd1 vccd1 vccd1 HI[74] insts\[74\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[207\] vssd1 vssd1 vccd1 vccd1 HI[207] insts\[207\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[157\] vssd1 vssd1 vccd1 vccd1 HI[157] insts\[157\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[324\] vssd1 vssd1 vccd1 vccd1 HI[324] insts\[324\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[37\] vssd1 vssd1 vccd1 vccd1 HI[37] insts\[37\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[441\] vssd1 vssd1 vccd1 vccd1 HI[441] insts\[441\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[274\] vssd1 vssd1 vccd1 vccd1 HI[274] insts\[274\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[391\] vssd1 vssd1 vccd1 vccd1 HI[391] insts\[391\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[237\] vssd1 vssd1 vccd1 vccd1 HI[237] insts\[237\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[404\] vssd1 vssd1 vccd1 vccd1 HI[404] insts\[404\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[354\] vssd1 vssd1 vccd1 vccd1 HI[354] insts\[354\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[187\] vssd1 vssd1 vccd1 vccd1 HI[187] insts\[187\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[67\] vssd1 vssd1 vccd1 vccd1 HI[67] insts\[67\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[102\] vssd1 vssd1 vccd1 vccd1 HI[102] insts\[102\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[317\] vssd1 vssd1 vccd1 vccd1 HI[317] insts\[317\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[434\] vssd1 vssd1 vccd1 vccd1 HI[434] insts\[434\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[267\] vssd1 vssd1 vccd1 vccd1 HI[267] insts\[267\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[384\] vssd1 vssd1 vccd1 vccd1 HI[384] insts\[384\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[97\] vssd1 vssd1 vccd1 vccd1 HI[97] insts\[97\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[132\] vssd1 vssd1 vccd1 vccd1 HI[132] insts\[132\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[12\] vssd1 vssd1 vccd1 vccd1 HI[12] insts\[12\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[347\] vssd1 vssd1 vccd1 vccd1 HI[347] insts\[347\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[297\] vssd1 vssd1 vccd1 vccd1 HI[297] insts\[297\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[212\] vssd1 vssd1 vccd1 vccd1 HI[212] insts\[212\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[162\] vssd1 vssd1 vccd1 vccd1 HI[162] insts\[162\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[427\] vssd1 vssd1 vccd1 vccd1 HI[427] insts\[427\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[42\] vssd1 vssd1 vccd1 vccd1 HI[42] insts\[42\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[377\] vssd1 vssd1 vccd1 vccd1 HI[377] insts\[377\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[0\] vssd1 vssd1 vccd1 vccd1 HI[0] insts\[0\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[125\] vssd1 vssd1 vccd1 vccd1 HI[125] insts\[125\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[242\] vssd1 vssd1 vccd1 vccd1 HI[242] insts\[242\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[457\] vssd1 vssd1 vccd1 vccd1 HI[457] insts\[457\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[192\] vssd1 vssd1 vccd1 vccd1 HI[192] insts\[192\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[72\] vssd1 vssd1 vccd1 vccd1 HI[72] insts\[72\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[205\] vssd1 vssd1 vccd1 vccd1 HI[205] insts\[205\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[155\] vssd1 vssd1 vccd1 vccd1 HI[155] insts\[155\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[322\] vssd1 vssd1 vccd1 vccd1 HI[322] insts\[322\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[35\] vssd1 vssd1 vccd1 vccd1 HI[35] insts\[35\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[272\] vssd1 vssd1 vccd1 vccd1 HI[272] insts\[272\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[118\] vssd1 vssd1 vccd1 vccd1 HI[118] insts\[118\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[235\] vssd1 vssd1 vccd1 vccd1 HI[235] insts\[235\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[402\] vssd1 vssd1 vccd1 vccd1 HI[402] insts\[402\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[185\] vssd1 vssd1 vccd1 vccd1 HI[185] insts\[185\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[352\] vssd1 vssd1 vccd1 vccd1 HI[352] insts\[352\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[65\] vssd1 vssd1 vccd1 vccd1 HI[65] insts\[65\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[100\] vssd1 vssd1 vccd1 vccd1 HI[100] insts\[100\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[148\] vssd1 vssd1 vccd1 vccd1 HI[148] insts\[148\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[315\] vssd1 vssd1 vccd1 vccd1 HI[315] insts\[315\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[28\] vssd1 vssd1 vccd1 vccd1 HI[28] insts\[28\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[265\] vssd1 vssd1 vccd1 vccd1 HI[265] insts\[265\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[432\] vssd1 vssd1 vccd1 vccd1 HI[432] insts\[432\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[382\] vssd1 vssd1 vccd1 vccd1 HI[382] insts\[382\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[95\] vssd1 vssd1 vccd1 vccd1 HI[95] insts\[95\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[228\] vssd1 vssd1 vccd1 vccd1 HI[228] insts\[228\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[130\] vssd1 vssd1 vccd1 vccd1 HI[130] insts\[130\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[10\] vssd1 vssd1 vccd1 vccd1 HI[10] insts\[10\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[178\] vssd1 vssd1 vccd1 vccd1 HI[178] insts\[178\]/LO sky130_fd_sc_hd__conb_1
XFILLER_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[345\] vssd1 vssd1 vccd1 vccd1 HI[345] insts\[345\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[58\] vssd1 vssd1 vccd1 vccd1 HI[58] insts\[58\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[295\] vssd1 vssd1 vccd1 vccd1 HI[295] insts\[295\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
.ends

.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
R0 VGND LO sky130_fd_pr__res_generic_po w=510000u l=45000u
R1 HI VPWR sky130_fd_pr__res_generic_po w=510000u l=45000u
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt mgmt_protect_hv vdda1 vssd vccd vdda2 mprj2_vdd_logic1 mprj_vdd_logic1
Xmprj2_logic_high_hvl vssd vssd vdda2 vdda2 mprj2_logic_high_lv/A mprj2_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_hvl vssd vssd vdda1 vdda1 mprj_logic_high_lv/A mprj_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_lv mprj_logic_high_lv/A vccd vssd vssd vdda1 vdda1 mprj_vdd_logic1
+ sky130_fd_sc_hvl__lsbufhv2lv_1
Xmprj2_logic_high_lv mprj2_logic_high_lv/A vccd vssd vssd vdda2 vdda2 mprj2_vdd_logic1
+ sky130_fd_sc_hvl__lsbufhv2lv_1
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12] mprj_adr_o_core[13]
+ mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16] mprj_adr_o_core[17]
+ mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21]
+ mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24] mprj_adr_o_core[25]
+ mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28] mprj_adr_o_core[29]
+ mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3] mprj_adr_o_core[4]
+ mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8] mprj_adr_o_core[9]
+ mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12] mprj_adr_o_user[13]
+ mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16] mprj_adr_o_user[17]
+ mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21]
+ mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24] mprj_adr_o_user[25]
+ mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28] mprj_adr_o_user[29]
+ mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3] mprj_adr_o_user[4]
+ mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8] mprj_adr_o_user[9]
+ mprj_cyc_o_core mprj_cyc_o_user mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11]
+ mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14] mprj_dat_o_core[15]
+ mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18] mprj_dat_o_core[19]
+ mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22] mprj_dat_o_core[23]
+ mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26] mprj_dat_o_core[27]
+ mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31]
+ mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7]
+ mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11]
+ mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14] mprj_dat_o_user[15]
+ mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18] mprj_dat_o_user[19]
+ mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22] mprj_dat_o_user[23]
+ mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26] mprj_dat_o_user[27]
+ mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31]
+ mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7]
+ mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2]
+ mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3]
+ mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood
+ user1_vdd_powergood user2_vcc_powergood user2_vdd_powergood user_clock user_clock2
+ user_irq[0] user_irq[1] user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2]
+ user_irq_ena[0] user_irq_ena[1] user_irq_ena[2] user_reset vccd vssd vccd1 vccd2
+ vdda1 vdda2
XFILLER_23_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[72\] la_iena_mprj[72] mprj_logic_high_inst/HI[402] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[72\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_501_ la_data_out_mprj[39] vssd vssd vccd vccd _501_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[50\] la_oenb_mprj[50] la_buf_enable\[50\]/B vssd vssd vccd vccd la_buf\[50\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_432_ mprj_dat_o_core[2] vssd vssd vccd vccd _432_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_363_ la_oenb_mprj[102] vssd vssd vccd vccd _363_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[36\] _498_/Y la_buf\[36\]/TE vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_35_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[108\] la_iena_mprj[108] mprj_logic_high_inst/HI[438] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[108\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] user_to_mprj_in_gates\[25\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[25\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_25_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[76\] _337_/Y mprj_logic_high_inst/HI[278] vssd vssd vccd
+ vccd la_oenb_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_26_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[98\] la_oenb_mprj[98] la_buf_enable\[98\]/B vssd vssd vccd vccd la_buf\[98\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[24\] _454_/Y mprj_dat_buf\[24\]/TE vssd vssd vccd vccd mprj_dat_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high_inst/HI[306] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_415_ mprj_adr_o_core[17] vssd vssd vccd vccd _415_/Y sky130_fd_sc_hd__inv_2
X_346_ la_oenb_mprj[85] vssd vssd vccd vccd _346_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[122\]_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[4\] la_oenb_mprj[4] la_buf_enable\[4\]/B vssd vssd vccd vccd la_buf\[4\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_9_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high_inst/HI[329] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[113\]_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[35\] la_iena_mprj[35] mprj_logic_high_inst/HI[365] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[35\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[13\] la_oenb_mprj[13] la_buf_enable\[13\]/B vssd vssd vccd vccd la_buf\[13\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[26\]_TE mprj_logic_high_inst/HI[228] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[92\]_A_N la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[104\]_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[30\]_A_N la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_329_ la_oenb_mprj[68] vssd vssd vccd vccd _329_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[45\]_A_N la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] user_to_mprj_in_gates\[92\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[92\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[64\]_TE la_buf\[64\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high_inst/HI[251] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[109\] _370_/Y mprj_logic_high_inst/HI[311] vssd vssd vccd
+ vccd la_oenb_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_1_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[93\]_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[39\] _629_/Y mprj_logic_high_inst/HI[241] vssd vssd vccd
+ vccd la_oenb_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_34_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[13\]_TE mprj_dat_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__402__A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[84\]_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y vssd vssd vccd vccd la_data_in_mprj[62]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[75\]_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[80\] la_oenb_mprj[80] la_buf_enable\[80\]/B vssd vssd vccd vccd la_buf\[80\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[66\]_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[66\] _528_/Y la_buf\[66\]/TE vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__einvp_8
X_594_ la_oenb_mprj[4] vssd vssd vccd vccd _594_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[122\] _584_/Y la_buf\[122\]/TE vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__einvp_8
XFILLER_6_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[57\]_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] user_to_mprj_in_gates\[55\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[55\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[48\]_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[39\]_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_646_ la_oenb_mprj[56] vssd vssd vccd vccd _646_/Y sky130_fd_sc_hd__inv_2
X_577_ la_data_out_mprj[115] vssd vssd vccd vccd _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[6\]_A _436_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y vssd vssd vccd vccd la_data_in_mprj[25]
+ sky130_fd_sc_hd__inv_8
XFILLER_10_1290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__500__A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[65\] la_iena_mprj[65] mprj_logic_high_inst/HI[395] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[65\]/B sky130_fd_sc_hd__and2_1
X_500_ la_data_out_mprj[38] vssd vssd vccd vccd _500_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[3\] _593_/Y mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd la_oenb_core[3] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[21\] _611_/Y mprj_logic_high_inst/HI[223] vssd vssd vccd
+ vccd la_oenb_core[21] sky130_fd_sc_hd__einvp_8
X_431_ mprj_dat_o_core[1] vssd vssd vccd vccd _431_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[43\] la_oenb_mprj[43] la_buf_enable\[43\]/B vssd vssd vccd vccd la_buf\[43\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_362_ la_oenb_mprj[101] vssd vssd vccd vccd _362_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[29\] _491_/Y la_buf\[29\]/TE vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_29_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__410__A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_629_ la_oenb_mprj[39] vssd vssd vccd vccd _629_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] user_to_mprj_in_gates\[18\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[18\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high_inst/HI[284] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[69\] _330_/Y mprj_logic_high_inst/HI[271] vssd vssd vccd
+ vccd la_oenb_core[69] sky130_fd_sc_hd__einvp_8
XFILLER_8_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[17\] _447_/Y mprj_dat_buf\[17\]/TE vssd vssd vccd vccd mprj_dat_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_414_ mprj_adr_o_core[16] vssd vssd vccd vccd _414_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_345_ la_oenb_mprj[84] vssd vssd vccd vccd _345_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[120\] la_iena_mprj[120] mprj_logic_high_inst/HI[450] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[120\]/B sky130_fd_sc_hd__and2_1
XFILLER_15_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__405__A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[12\] _410_/Y mprj_adr_buf\[12\]/TE vssd vssd vccd vccd mprj_adr_o_user[12]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[126] sky130_fd_sc_hd__inv_8
XANTENNA_la_buf_enable\[50\]_B la_buf_enable\[50\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y vssd vssd vccd vccd la_data_in_mprj[92]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[122\]_B mprj_logic_high_inst/HI[452] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_A _485_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[41\]_B la_buf_enable\[41\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[113\]_B mprj_logic_high_inst/HI[443] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[28\] la_iena_mprj[28] mprj_logic_high_inst/HI[358] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[28\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[14\]_A _476_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[32\]_B la_buf_enable\[32\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[1\]_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[96\] _558_/Y la_buf\[96\]/TE vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[1\] la_iena_mprj[1] mprj_logic_high_inst/HI[331] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[1\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[111\] la_oenb_mprj[111] la_buf_enable\[111\]/B vssd vssd vccd vccd
+ la_buf\[111\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[104\]_B mprj_logic_high_inst/HI[434] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[99\]_B la_buf_enable\[99\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[23\]_B la_buf_enable\[23\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] user_to_mprj_in_gates\[85\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[85\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[14\]_B la_buf_enable\[14\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[93\]_B mprj_logic_high_inst/HI[423] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[7\] _469_/Y la_buf\[7\]/TE vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__einvp_8
XFILLER_10_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[11\] _473_/Y la_buf\[11\]/TE vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__einvp_8
XFILLER_4_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[4\] _402_/Y mprj_adr_buf\[4\]/TE vssd vssd vccd vccd mprj_adr_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[84\]_B mprj_logic_high_inst/HI[414] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y vssd vssd vccd vccd la_data_in_mprj[55]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high_inst/HI[319] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[75\]_B mprj_logic_high_inst/HI[405] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] user_to_mprj_in_gates\[111\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[111\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high_inst/HI[218] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[91\]_A_N la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__503__A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[95\] la_iena_mprj[95] mprj_logic_high_inst/HI[425] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[95\]/B sky130_fd_sc_hd__and2_1
XFILLER_20_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[121\] _382_/Y mprj_logic_high_inst/HI[323] vssd vssd vccd
+ vccd la_oenb_core[121] sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[2\] _396_/Y mprj_sel_buf\[2\]/TE vssd vssd vccd vccd mprj_sel_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[66\]_B mprj_logic_high_inst/HI[396] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[51\] _641_/Y mprj_logic_high_inst/HI[253] vssd vssd vccd
+ vccd la_oenb_core[51] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[73\] la_oenb_mprj[73] la_buf_enable\[73\]/B vssd vssd vccd vccd la_buf\[73\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[44\]_A_N la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_593_ la_oenb_mprj[3] vssd vssd vccd vccd _593_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[59\] _521_/Y la_buf\[59\]/TE vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[59\]_A_N la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__413__A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[115\] _577_/Y la_buf\[115\]/TE vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_10_1472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[57\]_B mprj_logic_high_inst/HI[387] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[54\]_TE la_buf\[54\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[39\]_TE mprj_logic_high_inst/HI[241] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] user_to_mprj_in_gates\[48\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[48\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_34_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[48\]_B mprj_logic_high_inst/HI[378] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[10\] la_iena_mprj[10] mprj_logic_high_inst/HI[340] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[10\]/B sky130_fd_sc_hd__and2_1
XFILLER_21_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[99\] _360_/Y mprj_logic_high_inst/HI[301] vssd vssd vccd
+ vccd la_oenb_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_5_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_vdd_pwrgood mprj2_vdd_pwrgood/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_1_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[39\]_B mprj_logic_high_inst/HI[369] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_645_ la_oenb_mprj[55] vssd vssd vccd vccd _645_/Y sky130_fd_sc_hd__inv_2
X_576_ la_data_out_mprj[114] vssd vssd vccd vccd _576_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__408__A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y vssd vssd vccd vccd la_data_in_mprj[18]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_adr_buf\[25\]_A _423_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[5\]_TE mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_A _414_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[58\] la_iena_mprj[58] mprj_logic_high_inst/HI[388] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[58\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_430_ mprj_dat_o_core[0] vssd vssd vccd vccd _430_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[14\] _604_/Y mprj_logic_high_inst/HI[216] vssd vssd vccd
+ vccd la_oenb_core[14] sky130_fd_sc_hd__einvp_8
X_361_ la_oenb_mprj[100] vssd vssd vccd vccd _361_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[36\] la_oenb_mprj[36] la_buf_enable\[36\]/B vssd vssd vccd vccd la_buf\[36\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_628_ la_oenb_mprj[38] vssd vssd vccd vccd _628_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_559_ la_data_out_mprj[97] vssd vssd vccd vccd _559_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__601__A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__511__A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_413_ mprj_adr_o_core[15] vssd vssd vccd vccd _413_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[41\] _503_/Y la_buf\[41\]/TE vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[102\]_TE la_buf\[102\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_344_ la_oenb_mprj[83] vssd vssd vccd vccd _344_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[113\] la_iena_mprj[113] mprj_logic_high_inst/HI[443] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[113\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[17\]_TE mprj_adr_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__421__A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[119] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[29\]_A _459_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y vssd vssd vccd vccd la_data_in_mprj[85]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] user_to_mprj_in_gates\[30\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[30\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_470 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__331__A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__506__A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[81\] _342_/Y mprj_logic_high_inst/HI[283] vssd vssd vccd
+ vccd la_oenb_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_2_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[1\]_B mprj_logic_high_inst/HI[331] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[89\] _551_/Y la_buf\[89\]/TE vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_0_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[104\] la_oenb_mprj[104] la_buf_enable\[104\]/B vssd vssd vccd vccd
+ la_buf\[104\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_0_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[72\]_TE mprj_logic_high_inst/HI[274] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__416__A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] user_to_mprj_in_gates\[78\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[78\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[122\]_B la_buf_enable\[122\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[113\]_B la_buf_enable\[113\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[40\] la_iena_mprj[40] mprj_logic_high_inst/HI[370] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[40\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high_inst/HI[297] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[7\]_A _469_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[104\]_B la_buf_enable\[104\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y vssd vssd vccd vccd la_data_in_mprj[48]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] user_to_mprj_in_gates\[104\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[104\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[88\] la_iena_mprj[88] mprj_logic_high_inst/HI[418] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[88\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[114\] _375_/Y mprj_logic_high_inst/HI[316] vssd vssd vccd
+ vccd la_oenb_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_5_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[44\] _634_/Y mprj_logic_high_inst/HI[246] vssd vssd vccd
+ vccd la_oenb_core[44] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[66\] la_oenb_mprj[66] la_buf_enable\[66\]/B vssd vssd vccd vccd la_buf\[66\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_irq_buffers\[2\] user_irq_gates\[2\]/Y vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__inv_8
X_592_ la_oenb_mprj[2] vssd vssd vccd vccd _592_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[108\] _570_/Y la_buf\[108\]/TE vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__einvp_8
XFILLER_3_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[101] sky130_fd_sc_hd__inv_8
XFILLER_3_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__604__A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[0\] _430_/Y mprj_dat_buf\[0\]/TE vssd vssd vccd vccd mprj_dat_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__514__A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_644_ la_oenb_mprj[54] vssd vssd vccd vccd _644_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[71\] _533_/Y la_buf\[71\]/TE vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__einvp_8
X_575_ la_data_out_mprj[113] vssd vssd vccd vccd _575_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__424__A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[90\]_A_N la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] user_to_mprj_in_gates\[60\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[60\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__334__A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_30_1646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[43\]_A_N la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[58\]_A_N la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__509__A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_360_ la_oenb_mprj[99] vssd vssd vccd vccd _360_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[29\] la_oenb_mprj[29] la_buf_enable\[29\]/B vssd vssd vccd vccd la_buf\[29\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_10_810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high_inst/HI[231] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__419__A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_627_ la_oenb_mprj[37] vssd vssd vccd vccd _627_/Y sky130_fd_sc_hd__inv_2
X_558_ la_data_out_mprj[96] vssd vssd vccd vccd _558_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y vssd vssd vccd vccd la_data_in_mprj[30]
+ sky130_fd_sc_hd__inv_8
X_489_ la_data_out_mprj[27] vssd vssd vccd vccd _489_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[1\]_B la_buf_enable\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[125\]_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__329__A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[70\] la_iena_mprj[70] mprj_logic_high_inst/HI[400] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[70\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[116\]_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_412_ mprj_adr_o_core[14] vssd vssd vccd vccd _412_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_343_ la_oenb_mprj[82] vssd vssd vccd vccd _343_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[34\] _496_/Y la_buf\[34\]/TE vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[106\] la_iena_mprj[106] mprj_logic_high_inst/HI[436] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[106\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[107\]_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y vssd vssd vccd vccd la_data_in_mprj[78]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] user_to_mprj_in_gates\[23\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[23\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__612__A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__522__A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[74\] _335_/Y mprj_logic_high_inst/HI[276] vssd vssd vccd
+ vccd la_oenb_core[74] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[96\] la_oenb_mprj[96] la_buf_enable\[96\]/B vssd vssd vccd vccd la_buf\[96\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[96\]_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[22\] _452_/Y mprj_dat_buf\[22\]/TE vssd vssd vccd vccd mprj_dat_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[20\]_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__432__A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[87\]_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__607__A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[11\]_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[2\] la_oenb_mprj[2] la_buf_enable\[2\]/B vssd vssd vccd vccd la_buf\[2\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__342__A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[78\]_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[33\] la_iena_mprj[33] mprj_logic_high_inst/HI[363] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[33\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__517__A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[11\] la_oenb_mprj[11] la_buf_enable\[11\]/B vssd vssd vccd vccd la_buf\[11\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_3_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[69\]_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__427__A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] user_to_mprj_in_gates\[90\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[90\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__337__A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[62\]_TE mprj_logic_high_inst/HI[264] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[107\] _368_/Y mprj_logic_high_inst/HI[309] vssd vssd vccd
+ vccd la_oenb_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_5_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[37\] _627_/Y mprj_logic_high_inst/HI[239] vssd vssd vccd
+ vccd la_oenb_core[37] sky130_fd_sc_hd__einvp_8
X_591_ la_oenb_mprj[1] vssd vssd vccd vccd _591_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[59\] la_oenb_mprj[59] la_buf_enable\[59\]/B vssd vssd vccd vccd la_buf\[59\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y vssd vssd vccd vccd la_data_in_mprj[60]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[9\]_A _439_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[80\]_A _542_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high_inst/HI[287] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__620__A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[71\]_A _533_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__530__A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_643_ la_oenb_mprj[53] vssd vssd vccd vccd _643_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[64\] _526_/Y la_buf\[64\]/TE vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__einvp_8
X_574_ la_data_out_mprj[112] vssd vssd vccd vccd _574_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[62\]_A _524_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B user_to_mprj_in_gates\[112\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[28\] _426_/Y mprj_adr_buf\[28\]/TE vssd vssd vccd vccd mprj_adr_o_user[28]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[120\] _582_/Y la_buf\[120\]/TE vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[80\]_B la_buf_enable\[80\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__440__A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] user_to_mprj_in_gates\[53\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[53\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__615__A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[53\]_A _515_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[71\]_B la_buf_enable\[71\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__350__A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__525__A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[127\] la_oenb_mprj[127] la_buf_enable\[127\]/B vssd vssd vccd vccd
+ la_buf\[127\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_20_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_626_ la_oenb_mprj[36] vssd vssd vccd vccd _626_/Y sky130_fd_sc_hd__inv_2
X_557_ la_data_out_mprj[95] vssd vssd vccd vccd _557_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__435__A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_488_ la_data_out_mprj[26] vssd vssd vccd vccd _488_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y vssd vssd vccd vccd la_data_in_mprj[23]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf_enable\[53\]_B la_buf_enable\[53\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[125\]_B mprj_logic_high_inst/HI[455] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__345__A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_A _488_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[44\]_B la_buf_enable\[44\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[63\] la_iena_mprj[63] mprj_logic_high_inst/HI[393] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[63\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[116\]_B mprj_logic_high_inst/HI[446] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[1\] _591_/Y mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd la_oenb_core[1] sky130_fd_sc_hd__einvp_8
X_411_ mprj_adr_o_core[13] vssd vssd vccd vccd _411_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[41\] la_oenb_mprj[41] la_buf_enable\[41\]/B vssd vssd vccd vccd la_buf\[41\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_342_ la_oenb_mprj[81] vssd vssd vccd vccd _342_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[17\]_A _479_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[27\] _489_/Y la_buf\[27\]/TE vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__einvp_8
XFILLER_10_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[35\]_B la_buf_enable\[35\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[4\]_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[102\]_A _363_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[107\]_B mprj_logic_high_inst/HI[437] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[42\]_A_N la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_609_ la_oenb_mprj[19] vssd vssd vccd vccd _609_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] user_to_mprj_in_gates\[16\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[16\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[57\]_A_N la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[26\]_B la_buf_enable\[26\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] user_to_mprj_in_gates\[127\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[127\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[34\]_TE la_buf\[34\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high_inst/HI[221] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[17\]_B la_buf_enable\[17\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[96\]_B mprj_logic_high_inst/HI[426] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[67\] _657_/Y mprj_logic_high_inst/HI[269] vssd vssd vccd
+ vccd la_oenb_core[67] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[89\] la_oenb_mprj[89] la_buf_enable\[89\]/B vssd vssd vccd vccd la_buf\[89\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[15\] _445_/Y mprj_dat_buf\[15\]/TE vssd vssd vccd vccd mprj_dat_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_27_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[20\]_B mprj_logic_high_inst/HI[350] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[10\] _408_/Y mprj_adr_buf\[10\]/TE vssd vssd vccd vccd mprj_adr_o_user[10]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[124] sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[87\]_B mprj_logic_high_inst/HI[417] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y vssd vssd vccd vccd la_data_in_mprj[90]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[11\]_B mprj_logic_high_inst/HI[341] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__623__A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[26\] la_iena_mprj[26] mprj_logic_high_inst/HI[356] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[26\]/B sky130_fd_sc_hd__and2_1
XFILLER_32_1314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__533__A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[94\] _556_/Y la_buf\[94\]/TE vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_1_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__443__A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] user_to_mprj_in_gates\[83\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[83\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__618__A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__353__A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_590_ la_oenb_mprj[0] vssd vssd vccd vccd _590_/Y sky130_fd_sc_hd__inv_2
XANTENNA__528__A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[5\] _467_/Y la_buf\[5\]/TE vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__einvp_8
XFILLER_3_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[2\] _400_/Y mprj_adr_buf\[2\]/TE vssd vssd vccd vccd mprj_adr_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_35_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__438__A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y vssd vssd vccd vccd la_data_in_mprj[53]
+ sky130_fd_sc_hd__inv_8
XFILLER_35_658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[28\]_A _426_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__348__A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[93\] la_iena_mprj[93] mprj_logic_high_inst/HI[423] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[93\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_sel_buf\[0\] _394_/Y mprj_sel_buf\[0\]/TE vssd vssd vccd vccd mprj_sel_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[71\] la_oenb_mprj[71] la_buf_enable\[71\]/B vssd vssd vccd vccd la_buf\[71\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_642_ la_oenb_mprj[52] vssd vssd vccd vccd _642_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_573_ la_data_out_mprj[111] vssd vssd vccd vccd _573_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[57\] _519_/Y la_buf\[57\]/TE vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__einvp_8
XFILLER_18_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[113\] _575_/Y la_buf\[113\]/TE vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__einvp_8
XFILLER_23_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] user_to_mprj_in_gates\[46\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[46\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high_inst/HI[254] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__631__A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] user_to_mprj_in_gates\[8\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[8\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[97\] _358_/Y mprj_logic_high_inst/HI[299] vssd vssd vccd
+ vccd la_oenb_core[97] sky130_fd_sc_hd__einvp_8
XFILLER_5_348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__541__A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_625_ la_oenb_mprj[35] vssd vssd vccd vccd _625_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high_inst/HI[277] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_556_ la_data_out_mprj[94] vssd vssd vccd vccd _556_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_487_ la_data_out_mprj[25] vssd vssd vccd vccd _487_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y vssd vssd vccd vccd la_data_in_mprj[16]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__451__A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__626__A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[4\]_A _402_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__361__A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[56\] la_iena_mprj[56] mprj_logic_high_inst/HI[386] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[56\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high_inst/HI[300] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_410_ mprj_adr_o_core[12] vssd vssd vccd vccd _410_/Y sky130_fd_sc_hd__inv_2
XANTENNA__536__A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[12\] _602_/Y mprj_logic_high_inst/HI[214] vssd vssd vccd
+ vccd la_oenb_core[12] sky130_fd_sc_hd__einvp_8
X_341_ la_oenb_mprj[80] vssd vssd vccd vccd _341_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[34\] la_oenb_mprj[34] la_buf_enable\[34\]/B vssd vssd vccd vccd la_buf\[34\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y vssd vssd vccd vccd la_data_in_mprj[8]
+ sky130_fd_sc_hd__inv_8
XFILLER_17_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[4\]_B mprj_logic_high_inst/HI[334] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_stb_buf _392_/Y mprj_stb_buf/TE vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__einvp_8
XFILLER_2_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_608_ la_oenb_mprj[18] vssd vssd vccd vccd _608_/Y sky130_fd_sc_hd__inv_2
XANTENNA__446__A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_539_ la_data_out_mprj[77] vssd vssd vccd vccd _539_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[125\]_B la_buf_enable\[125\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__356__A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[116\]_B la_buf_enable\[116\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[111\] la_iena_mprj[111] mprj_logic_high_inst/HI[441] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[111\]/B sky130_fd_sc_hd__and2_1
XFILLER_7_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[30\]_TE mprj_adr_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[117] sky130_fd_sc_hd__inv_8
XFILLER_6_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y vssd vssd vccd vccd la_data_in_mprj[83]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf_enable\[107\]_B la_buf_enable\[107\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[19\] la_iena_mprj[19] mprj_logic_high_inst/HI[349] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[19\]/B sky130_fd_sc_hd__and2_1
XFILLER_32_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[41\]_A_N la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[56\]_A_N la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[87\] _549_/Y la_buf\[87\]/TE vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_21_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[102\] la_oenb_mprj[102] la_buf_enable\[102\]/B vssd vssd vccd vccd
+ la_buf\[102\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_1_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_TE la_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] user_to_mprj_in_gates\[76\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[76\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__634__A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2050 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_2083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__544__A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_ena_buf\[2\] user_irq_ena[2] user_irq_ena_buf\[2\]/B vssd vssd vccd vccd
+ user_irq_gates\[2\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y vssd vssd vccd vccd la_data_in_mprj[46]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__454__A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__629__A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] user_to_mprj_in_gates\[102\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[102\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__364__A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[86\] la_iena_mprj[86] mprj_logic_high_inst/HI[416] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[86\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[112\] _373_/Y mprj_logic_high_inst/HI[314] vssd vssd vccd
+ vccd la_oenb_core[112] sky130_fd_sc_hd__einvp_8
XANTENNA__539__A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[42\] _632_/Y mprj_logic_high_inst/HI[244] vssd vssd vccd
+ vccd la_oenb_core[42] sky130_fd_sc_hd__einvp_8
X_641_ la_oenb_mprj[51] vssd vssd vccd vccd _641_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[64\] la_oenb_mprj[64] la_buf_enable\[64\]/B vssd vssd vccd vccd la_buf\[64\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_irq_buffers\[0\] user_irq_gates\[0\]/Y vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__inv_8
X_572_ la_data_out_mprj[110] vssd vssd vccd vccd _572_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[106\] _568_/Y la_buf\[106\]/TE vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__einvp_8
XFILLER_7_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__449__A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] user_to_mprj_in_gates\[39\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[39\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1059 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[4\]_B la_buf_enable\[4\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__359__A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[119\]_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high_inst/HI[322] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_624_ la_oenb_mprj[34] vssd vssd vccd vccd _624_/Y sky130_fd_sc_hd__inv_2
X_555_ la_data_out_mprj[93] vssd vssd vccd vccd _555_/Y sky130_fd_sc_hd__inv_2
X_486_ la_data_out_mprj[24] vssd vssd vccd vccd _486_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[50\]_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_we_buf _393_/Y mprj_we_buf/TE vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__einvp_8
XFILLER_9_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_pwrgood mprj_pwrgood/A vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_9_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[41\]_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__642__A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[49\] la_iena_mprj[49] mprj_logic_high_inst/HI[379] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[49\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_340_ la_oenb_mprj[79] vssd vssd vccd vccd _340_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[32\]_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[27\] la_oenb_mprj[27] la_buf_enable\[27\]/B vssd vssd vccd vccd la_buf\[27\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__552__A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[99\]_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_607_ la_oenb_mprj[17] vssd vssd vccd vccd _607_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[23\]_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_538_ la_data_out_mprj[76] vssd vssd vccd vccd _538_/Y sky130_fd_sc_hd__inv_2
X_469_ la_data_out_mprj[7] vssd vssd vccd vccd _469_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__462__A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__637__A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[14\]_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__372__A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[65\]_TE mprj_logic_high_inst/HI[267] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1299 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__547__A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_ena_buf\[1\]_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_we_buf_A _393_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[32\] _494_/Y la_buf\[32\]/TE vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[104\] la_iena_mprj[104] mprj_logic_high_inst/HI[434] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[104\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y vssd vssd vccd vccd la_data_in_mprj[76]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__457__A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] user_to_mprj_in_gates\[21\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[21\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high_inst/HI[290] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[9\] _439_/Y mprj_dat_buf\[9\]/TE vssd vssd vccd vccd mprj_dat_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_2182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__367__A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[72\] _333_/Y mprj_logic_high_inst/HI[274] vssd vssd vccd
+ vccd la_oenb_core[72] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[94\] la_oenb_mprj[94] la_buf_enable\[94\]/B vssd vssd vccd vccd la_buf\[94\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[20\] _450_/Y mprj_dat_buf\[20\]/TE vssd vssd vccd vccd mprj_dat_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[92\]_A _554_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] user_to_mprj_in_gates\[69\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[69\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[83\]_A _545_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[0\] la_oenb_mprj[0] la_buf_enable\[0\]/B vssd vssd vccd vccd la_buf\[0\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__650__A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[31\] la_iena_mprj[31] mprj_logic_high_inst/HI[361] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[31\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[20\]_TE mprj_adr_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[74\]_A _536_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[124\]_B user_to_mprj_in_gates\[124\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[92\]_B la_buf_enable\[92\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__560__A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y vssd vssd vccd vccd la_data_in_mprj[39]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[65\]_A _527_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[83\]_B la_buf_enable\[83\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__470__A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__645__A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[40\]_A_N la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[106\]_B user_to_mprj_in_gates\[106\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[74\]_B la_buf_enable\[74\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[55\]_A_N la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__380__A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[79\] la_iena_mprj[79] mprj_logic_high_inst/HI[409] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[79\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[105\] _366_/Y mprj_logic_high_inst/HI[307] vssd vssd vccd
+ vccd la_oenb_core[105] sky130_fd_sc_hd__einvp_8
XFILLER_5_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_640_ la_oenb_mprj[50] vssd vssd vccd vccd _640_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[35\] _625_/Y mprj_logic_high_inst/HI[237] vssd vssd vccd
+ vccd la_oenb_core[35] sky130_fd_sc_hd__einvp_8
X_571_ la_data_out_mprj[109] vssd vssd vccd vccd _571_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[57\] la_oenb_mprj[57] la_buf_enable\[57\]/B vssd vssd vccd vccd la_buf\[57\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__555__A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[65\]_B la_buf_enable\[65\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__465__A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[56\]_B la_buf_enable\[56\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__375__A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[119\]_B mprj_logic_high_inst/HI[449] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_623_ la_oenb_mprj[33] vssd vssd vccd vccd _623_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[62\] _524_/Y la_buf\[62\]/TE vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__einvp_8
X_554_ la_data_out_mprj[92] vssd vssd vccd vccd _554_/Y sky130_fd_sc_hd__inv_2
X_485_ la_data_out_mprj[23] vssd vssd vccd vccd _485_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[50\]_B mprj_logic_high_inst/HI[380] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[38\]_B la_buf_enable\[38\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[7\]_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[26\] _424_/Y mprj_adr_buf\[26\]/TE vssd vssd vccd vccd mprj_adr_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] user_to_mprj_in_gates\[51\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[51\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[41\]_B mprj_logic_high_inst/HI[371] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[29\]_B la_buf_enable\[29\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[31\]_A _621_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[32\]_B mprj_logic_high_inst/HI[362] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[99\]_B mprj_logic_high_inst/HI[429] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[125\] la_oenb_mprj[125] la_buf_enable\[125\]/B vssd vssd vccd vccd
+ la_buf\[125\]/TE sky130_fd_sc_hd__and2b_1
X_606_ la_oenb_mprj[16] vssd vssd vccd vccd _606_/Y sky130_fd_sc_hd__inv_2
X_537_ la_data_out_mprj[75] vssd vssd vccd vccd _537_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[23\]_B mprj_logic_high_inst/HI[353] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_468_ la_data_out_mprj[6] vssd vssd vccd vccd _468_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_399_ mprj_adr_o_core[1] vssd vssd vccd vccd _399_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y vssd vssd vccd vccd la_data_in_mprj[21]
+ sky130_fd_sc_hd__inv_8
XFILLER_31_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] user_to_mprj_in_gates\[99\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[99\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[14\]_B mprj_logic_high_inst/HI[344] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__653__A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[110\]_TE mprj_logic_high_inst/HI[312] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[61\] la_iena_mprj[61] mprj_logic_high_inst/HI[391] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[61\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_ena_buf\[1\]_B user_irq_ena_buf\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__563__A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[25\] _487_/Y la_buf\[25\]/TE vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__einvp_8
XFILLER_1_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y vssd vssd vccd vccd la_data_in_mprj[69]
+ sky130_fd_sc_hd__inv_8
XANTENNA__473__A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] user_to_mprj_in_gates\[14\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[14\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] user_to_mprj_in_gates\[125\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[125\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__648__A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[31\]_A _461_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__383__A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[65\] _655_/Y mprj_logic_high_inst/HI[267] vssd vssd vccd
+ vccd la_oenb_core[65] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[87\] la_oenb_mprj[87] la_buf_enable\[87\]/B vssd vssd vccd vccd la_buf\[87\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[13\] _443_/Y mprj_dat_buf\[13\]/TE vssd vssd vccd vccd mprj_dat_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__558__A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[7\]_TE mprj_adr_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[122] sky130_fd_sc_hd__inv_8
XANTENNA__468__A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[13\]_A _443_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[55\]_TE mprj_logic_high_inst/HI[257] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__378__A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[24\] la_iena_mprj[24] mprj_logic_high_inst/HI[354] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[24\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[92\] _554_/Y la_buf\[92\]/TE vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_23_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high_inst/HI[280] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_31_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] user_to_mprj_in_gates\[81\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[81\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[9\]_A_N la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_570_ la_data_out_mprj[108] vssd vssd vccd vccd _570_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[28\] _618_/Y mprj_logic_high_inst/HI[230] vssd vssd vccd
+ vccd la_oenb_core[28] sky130_fd_sc_hd__einvp_8
XFILLER_12_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__571__A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[3\] _465_/Y la_buf\[3\]/TE vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__einvp_8
XFILLER_4_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[0\] _398_/Y mprj_adr_buf\[0\]/TE vssd vssd vccd vccd mprj_adr_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y vssd vssd vccd vccd la_data_in_mprj[51]
+ sky130_fd_sc_hd__inv_8
XFILLER_31_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__481__A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__656__A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[7\]_A _405_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__391__A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[91\] la_iena_mprj[91] mprj_logic_high_inst/HI[421] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[91\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_622_ la_oenb_mprj[32] vssd vssd vccd vccd _622_/Y sky130_fd_sc_hd__inv_2
XANTENNA__566__A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_553_ la_data_out_mprj[91] vssd vssd vccd vccd _553_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[55\] _517_/Y la_buf\[55\]/TE vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__einvp_8
X_484_ la_data_out_mprj[22] vssd vssd vccd vccd _484_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[127\] la_iena_mprj[127] mprj_logic_high_inst/HI[457] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[127\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[7\]_B mprj_logic_high_inst/HI[337] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[19\] _417_/Y mprj_adr_buf\[19\]/TE vssd vssd vccd vccd mprj_adr_o_user[19]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[111\] _573_/Y la_buf\[111\]/TE vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__einvp_8
XFILLER_4_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1083 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y vssd vssd vccd vccd la_data_in_mprj[99]
+ sky130_fd_sc_hd__inv_8
XFILLER_27_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[54\]_A_N la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__476__A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] user_to_mprj_in_gates\[44\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[44\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[69\]_A_N la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] user_to_mprj_in_gates\[6\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[6\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__386__A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[95\] _356_/Y mprj_logic_high_inst/HI[297] vssd vssd vccd
+ vccd la_oenb_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_5_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[119\]_B la_buf_enable\[119\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[8\] la_iena_mprj[8] mprj_logic_high_inst/HI[338] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[8\]/B sky130_fd_sc_hd__and2_1
XFILLER_37_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[118\] la_oenb_mprj[118] la_buf_enable\[118\]/B vssd vssd vccd vccd
+ la_buf\[118\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_605_ la_oenb_mprj[15] vssd vssd vccd vccd _605_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_536_ la_data_out_mprj[74] vssd vssd vccd vccd _536_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_467_ la_data_out_mprj[5] vssd vssd vccd vccd _467_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_398_ mprj_adr_o_core[0] vssd vssd vccd vccd _398_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y vssd vssd vccd vccd la_data_in_mprj[14]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[27\]_TE la_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[54\] la_iena_mprj[54] mprj_logic_high_inst/HI[384] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[54\]/B sky130_fd_sc_hd__and2_1
XFILLER_21_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[10\] _600_/Y mprj_logic_high_inst/HI[212] vssd vssd vccd
+ vccd la_oenb_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_19_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y vssd vssd vccd vccd la_data_in_mprj[6]
+ sky130_fd_sc_hd__inv_8
Xla_buf_enable\[32\] la_oenb_mprj[32] la_buf_enable\[32\]/B vssd vssd vccd vccd la_buf\[32\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[18\] _480_/Y la_buf\[18\]/TE vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_26_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_519_ la_data_out_mprj[57] vssd vssd vccd vccd _519_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_2223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] user_to_mprj_in_gates\[118\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[118\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[58\] _648_/Y mprj_logic_high_inst/HI[260] vssd vssd vccd
+ vccd la_oenb_core[58] sky130_fd_sc_hd__einvp_8
XFILLER_8_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__574__A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[100\]_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[115] sky130_fd_sc_hd__inv_8
XFILLER_26_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y vssd vssd vccd vccd la_data_in_mprj[81]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high_inst/HI[302] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__484__A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__394__A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_12_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[17\] la_iena_mprj[17] mprj_logic_high_inst/HI[347] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[17\]/B sky130_fd_sc_hd__and2_1
XFILLER_16_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__569__A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high_inst/HI[325] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[85\] _547_/Y la_buf\[85\]/TE vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_19_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[100\] la_oenb_mprj[100] la_buf_enable\[100\]/B vssd vssd vccd vccd
+ la_buf\[100\]/TE sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[80\]_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] user_to_mprj_in_gates\[74\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[74\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__479__A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[71\]_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[7\]_B la_buf_enable\[7\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__389__A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[62\]_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_ena_buf\[0\] user_irq_ena[0] user_irq_ena_buf\[0\]/B vssd vssd vccd vccd
+ user_irq_gates\[0\]/B sky130_fd_sc_hd__and2_1
XFILLER_7_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[53\]_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y vssd vssd vccd vccd la_data_in_mprj[44]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] user_to_mprj_in_gates\[100\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[100\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[44\]_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[84\] la_iena_mprj[84] mprj_logic_high_inst/HI[414] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[84\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[110\] _371_/Y mprj_logic_high_inst/HI[312] vssd vssd vccd
+ vccd la_oenb_core[110] sky130_fd_sc_hd__einvp_8
XFILLER_7_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[40\] _630_/Y mprj_logic_high_inst/HI[242] vssd vssd vccd
+ vccd la_oenb_core[40] sky130_fd_sc_hd__einvp_8
X_621_ la_oenb_mprj[31] vssd vssd vccd vccd _621_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[62\] la_oenb_mprj[62] la_buf_enable\[62\]/B vssd vssd vccd vccd la_buf\[62\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[35\]_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_552_ la_data_out_mprj[90] vssd vssd vccd vccd _552_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_483_ la_data_out_mprj[21] vssd vssd vccd vccd _483_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__582__A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[48\] _510_/Y la_buf\[48\]/TE vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_13_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[2\]_A _432_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[104\] _566_/Y la_buf\[104\]/TE vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_4_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[26\]_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] user_to_mprj_in_gates\[37\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[37\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__492__A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[8\]_A_N la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[17\]_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1382 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[88\] _349_/Y mprj_logic_high_inst/HI[290] vssd vssd vccd
+ vccd la_oenb_core[88] sky130_fd_sc_hd__einvp_8
XFILLER_1_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__577__A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_604_ la_oenb_mprj[14] vssd vssd vccd vccd _604_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_535_ la_data_out_mprj[73] vssd vssd vccd vccd _535_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_466_ la_data_out_mprj[4] vssd vssd vccd vccd _466_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_397_ mprj_sel_o_core[3] vssd vssd vccd vccd _397_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[31\] _429_/Y mprj_adr_buf\[31\]/TE vssd vssd vccd vccd mprj_adr_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_31_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__487__A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[100\]_A _562_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__397__A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[47\] la_iena_mprj[47] mprj_logic_high_inst/HI[377] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[47\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[23\]_TE mprj_adr_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[25\] la_oenb_mprj[25] la_buf_enable\[25\]/B vssd vssd vccd vccd la_buf\[25\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[53\]_A_N la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[68\]_A_N la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_A _557_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_518_ la_data_out_mprj[56] vssd vssd vccd vccd _518_/Y sky130_fd_sc_hd__inv_2
X_449_ mprj_dat_o_core[19] vssd vssd vccd vccd _449_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[86\]_A _548_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[10\]_A _472_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[100\]_B mprj_logic_high_inst/HI[430] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[95\]_B la_buf_enable\[95\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__590__A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[30\] _492_/Y la_buf\[30\]/TE vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[102\] la_iena_mprj[102] mprj_logic_high_inst/HI[432] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[102\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[108] sky130_fd_sc_hd__inv_8
XFILLER_6_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y vssd vssd vccd vccd la_data_in_mprj[74]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[118\]_B user_to_mprj_in_gates\[118\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[86\]_B la_buf_enable\[86\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[7\] _437_/Y mprj_dat_buf\[7\]/TE vssd vssd vccd vccd mprj_dat_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_2054 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[10\]_B la_buf_enable\[10\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[77\]_B la_buf_enable\[77\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[70\] _331_/Y mprj_logic_high_inst/HI[272] vssd vssd vccd
+ vccd la_oenb_core[70] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[92\] la_oenb_mprj[92] la_buf_enable\[92\]/B vssd vssd vccd vccd la_buf\[92\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[78\] _540_/Y la_buf\[78\]/TE vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__einvp_8
XFILLER_19_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__585__A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] user_to_mprj_in_gates\[67\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[67\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__495__A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[62\]_B mprj_logic_high_inst/HI[392] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[53\]_B mprj_logic_high_inst/HI[383] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y vssd vssd vccd vccd la_data_in_mprj[37]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[44\]_B mprj_logic_high_inst/HI[374] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high_inst/HI[315] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[77\] la_iena_mprj[77] mprj_logic_high_inst/HI[407] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[77\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[103\] _364_/Y mprj_logic_high_inst/HI[305] vssd vssd vccd
+ vccd la_oenb_core[103] sky130_fd_sc_hd__einvp_8
XFILLER_22_2361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_620_ la_oenb_mprj[30] vssd vssd vccd vccd _620_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[30\]_A _428_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[33\] _623_/Y mprj_logic_high_inst/HI[235] vssd vssd vccd
+ vccd la_oenb_core[33] sky130_fd_sc_hd__einvp_8
X_551_ la_data_out_mprj[89] vssd vssd vccd vccd _551_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[35\]_B mprj_logic_high_inst/HI[365] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[55\] la_oenb_mprj[55] la_buf_enable\[55\]/B vssd vssd vccd vccd la_buf\[55\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_482_ la_data_out_mprj[20] vssd vssd vccd vccd _482_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high_inst/HI[214] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_A _419_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[26\]_B mprj_logic_high_inst/HI[356] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_32_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[12\]_A _410_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[17\]_B mprj_logic_high_inst/HI[347] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high_inst/HI[237] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[109\]_A_N la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[29\] _459_/Y mprj_dat_buf\[29\]/TE vssd vssd vccd vccd mprj_dat_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_603_ la_oenb_mprj[13] vssd vssd vccd vccd _603_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[60\] _522_/Y la_buf\[60\]/TE vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__einvp_8
X_534_ la_data_out_mprj[72] vssd vssd vccd vccd _534_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__593__A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_465_ la_data_out_mprj[3] vssd vssd vccd vccd _465_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_396_ mprj_sel_o_core[2] vssd vssd vccd vccd _396_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[24\] _422_/Y mprj_adr_buf\[24\]/TE vssd vssd vccd vccd mprj_adr_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2005 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[9\] la_oenb_mprj[9] la_buf_enable\[9\]/B vssd vssd vccd vccd la_buf\[9\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_3_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[18\] la_oenb_mprj[18] la_buf_enable\[18\]/B vssd vssd vccd vccd la_buf\[18\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[1\]_TE mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_irq_gates\[1\] user_irq_core[1] user_irq_gates\[1\]/B vssd vssd vccd vccd user_irq_gates\[1\]/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_2_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__588__A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf_enable\[123\] la_oenb_mprj[123] la_buf_enable\[123\]/B vssd vssd vccd vccd
+ la_buf\[123\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_8_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[7\]_A_N la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[25\]_A _455_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_517_ la_data_out_mprj[55] vssd vssd vccd vccd _517_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_448_ mprj_dat_o_core[18] vssd vssd vccd vccd _448_/Y sky130_fd_sc_hd__inv_2
X_379_ la_oenb_mprj[118] vssd vssd vccd vccd _379_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] user_to_mprj_in_gates\[97\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[97\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__498__A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[16\]_A _446_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[23\] _485_/Y la_buf\[23\]/TE vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__einvp_8
XFILLER_10_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y vssd vssd vccd vccd la_data_in_mprj[67]
+ sky130_fd_sc_hd__inv_8
XFILLER_33_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] user_to_mprj_in_gates\[12\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[12\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[13\]_TE mprj_adr_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] user_to_mprj_in_gates\[123\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[123\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[52\]_A_N la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_A_N la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[63\] _653_/Y mprj_logic_high_inst/HI[265] vssd vssd vccd
+ vccd la_oenb_core[63] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[85\] la_oenb_mprj[85] la_buf_enable\[85\]/B vssd vssd vccd vccd la_buf\[85\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[11\] _441_/Y mprj_dat_buf\[11\]/TE vssd vssd vccd vccd mprj_dat_o_user[11]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_B la_buf_enable\[100\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[127\] _589_/Y la_buf\[127\]/TE vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__einvp_8
XFILLER_32_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[120] sky130_fd_sc_hd__inv_8
XFILLER_3_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[22\] la_iena_mprj[22] mprj_logic_high_inst/HI[352] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[22\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__596__A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[90\] _552_/Y la_buf\[90\]/TE vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_1_2158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high_inst/HI[293] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2071 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_550_ la_data_out_mprj[88] vssd vssd vccd vccd _550_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[26\] _616_/Y mprj_logic_high_inst/HI[228] vssd vssd vccd
+ vccd la_oenb_core[26] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[8\] _598_/Y mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd la_oenb_core[8] sky130_fd_sc_hd__einvp_8
X_481_ la_data_out_mprj[19] vssd vssd vccd vccd _481_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[48\] la_oenb_mprj[48] la_buf_enable\[48\]/B vssd vssd vccd vccd la_buf\[48\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[1\] _463_/Y la_buf\[1\]/TE vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_602_ la_oenb_mprj[12] vssd vssd vccd vccd _602_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_533_ la_data_out_mprj[71] vssd vssd vccd vccd _533_/Y sky130_fd_sc_hd__inv_2
X_464_ la_data_out_mprj[2] vssd vssd vccd vccd _464_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[53\] _515_/Y la_buf\[53\]/TE vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[125\] la_iena_mprj[125] mprj_logic_high_inst/HI[455] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[125\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_395_ mprj_sel_o_core[1] vssd vssd vccd vccd _395_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[17\] _415_/Y mprj_adr_buf\[17\]/TE vssd vssd vccd vccd mprj_adr_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y vssd vssd vccd vccd la_data_in_mprj[97]
+ sky130_fd_sc_hd__inv_8
XFILLER_29_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high_inst/HI[305] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] user_to_mprj_in_gates\[42\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[42\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[121\]_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] user_to_mprj_in_gates\[4\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[4\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[112\]_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[93\] _354_/Y mprj_logic_high_inst/HI[295] vssd vssd vccd
+ vccd la_oenb_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_2_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high_inst/HI[328] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[6\] la_iena_mprj[6] mprj_logic_high_inst/HI[336] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[6\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[116\] la_oenb_mprj[116] la_buf_enable\[116\]/B vssd vssd vccd vccd
+ la_buf\[116\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_2_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[103\]_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_516_ la_data_out_mprj[54] vssd vssd vccd vccd _516_/Y sky130_fd_sc_hd__inv_2
X_447_ mprj_dat_o_core[17] vssd vssd vccd vccd _447_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_378_ la_oenb_mprj[117] vssd vssd vccd vccd _378_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y vssd vssd vccd vccd la_data_in_mprj[12]
+ sky130_fd_sc_hd__inv_8
XFILLER_29_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[108\]_A_N la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[52\] la_iena_mprj[52] mprj_logic_high_inst/HI[382] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[52\]/B sky130_fd_sc_hd__and2_1
XFILLER_25_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[92\]_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y vssd vssd vccd vccd la_data_in_mprj[4]
+ sky130_fd_sc_hd__inv_8
Xla_buf_enable\[30\] la_oenb_mprj[30] la_buf_enable\[30\]/B vssd vssd vccd vccd la_buf\[30\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[16\] _478_/Y la_buf\[16\]/TE vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__einvp_8
XFILLER_10_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[48\]_TE mprj_logic_high_inst/HI[250] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__599__A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[9\] _407_/Y mprj_adr_buf\[9\]/TE vssd vssd vccd vccd mprj_adr_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[83\]_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] user_to_mprj_in_gates\[116\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[116\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[74\]_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[6\]_A_N la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[126\] _387_/Y mprj_logic_high_inst/HI[328] vssd vssd vccd
+ vccd la_oenb_core[126] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[56\] _646_/Y mprj_logic_high_inst/HI[258] vssd vssd vccd
+ vccd la_oenb_core[56] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[78\] la_oenb_mprj[78] la_buf_enable\[78\]/B vssd vssd vccd vccd la_buf\[78\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[65\]_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[113] sky130_fd_sc_hd__inv_8
XFILLER_3_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[56\]_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[47\]_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[15\] la_iena_mprj[15] mprj_logic_high_inst/HI[345] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[15\]/B sky130_fd_sc_hd__and2_1
XFILLER_21_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[38\]_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[83\] _545_/Y la_buf\[83\]/TE vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__einvp_8
XFILLER_5_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[5\]_A _435_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[51\]_A_N la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] user_to_mprj_in_gates\[72\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[72\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[66\]_A_N la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[29\]_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[19\]_A_N la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_480_ la_data_out_mprj[18] vssd vssd vccd vccd _480_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[19\] _609_/Y mprj_logic_high_inst/HI[221] vssd vssd vccd
+ vccd la_oenb_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_13_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__400__A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y vssd vssd vccd vccd la_data_in_mprj[42]
+ sky130_fd_sc_hd__inv_8
XFILLER_32_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[40\]_A _502_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[82\] la_iena_mprj[82] mprj_logic_high_inst/HI[412] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[82\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high_inst/HI[283] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_601_ la_oenb_mprj[11] vssd vssd vccd vccd _601_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[60\] la_oenb_mprj[60] la_buf_enable\[60\]/B vssd vssd vccd vccd la_buf\[60\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_532_ la_data_out_mprj[70] vssd vssd vccd vccd _532_/Y sky130_fd_sc_hd__inv_2
X_463_ la_data_out_mprj[1] vssd vssd vccd vccd _463_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[46\] _508_/Y la_buf\[46\]/TE vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__einvp_8
X_394_ mprj_sel_o_core[0] vssd vssd vccd vccd _394_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[118\] la_iena_mprj[118] mprj_logic_high_inst/HI[448] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[118\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[58\]_A user_to_mprj_in_gates\[58\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[102\] _564_/Y la_buf\[102\]/TE vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_7_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[121\]_B mprj_logic_high_inst/HI[451] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] user_to_mprj_in_gates\[35\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[35\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[22\]_A _484_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[40\]_B la_buf_enable\[40\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[89\]_A _551_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[112\]_B mprj_logic_high_inst/HI[442] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[13\]_A _475_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[86\] _347_/Y mprj_logic_high_inst/HI[288] vssd vssd vccd
+ vccd la_oenb_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_2_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[31\]_B la_buf_enable\[31\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[0\]_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[109\] la_oenb_mprj[109] la_buf_enable\[109\]/B vssd vssd vccd vccd
+ la_buf\[109\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_2_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[103\]_B mprj_logic_high_inst/HI[433] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_515_ la_data_out_mprj[53] vssd vssd vccd vccd _515_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[98\]_B la_buf_enable\[98\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_446_ mprj_dat_o_core[16] vssd vssd vccd vccd _446_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_377_ la_oenb_mprj[116] vssd vssd vccd vccd _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_B la_buf_enable\[22\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[89\]_B la_buf_enable\[89\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[13\]_B la_buf_enable\[13\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[92\]_B mprj_logic_high_inst/HI[422] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[45\] la_iena_mprj[45] mprj_logic_high_inst/HI[375] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[45\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[23\] la_oenb_mprj[23] la_buf_enable\[23\]/B vssd vssd vccd vccd la_buf\[23\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_23_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_429_ mprj_adr_o_core[31] vssd vssd vccd vccd _429_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] user_to_mprj_in_gates\[109\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[109\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high_inst/HI[318] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[119\] _380_/Y mprj_logic_high_inst/HI[321] vssd vssd vccd
+ vccd la_oenb_core[119] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[65\]_B mprj_logic_high_inst/HI[395] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[49\] _639_/Y mprj_logic_high_inst/HI[251] vssd vssd vccd
+ vccd la_oenb_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_15_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high_inst/HI[217] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[100\] la_iena_mprj[100] mprj_logic_high_inst/HI[430] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[100\]/B sky130_fd_sc_hd__and2_1
XANTENNA__403__A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[107\]_A_N la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[106] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y vssd vssd vccd vccd la_data_in_mprj[72]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[56\]_B mprj_logic_high_inst/HI[386] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[5\] _435_/Y mprj_dat_buf\[5\]/TE vssd vssd vccd vccd mprj_dat_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[47\]_B mprj_logic_high_inst/HI[377] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1855 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[38\]_TE mprj_logic_high_inst/HI[240] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[37\]_A _627_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[90\] la_oenb_mprj[90] la_buf_enable\[90\]/B vssd vssd vccd vccd la_buf\[90\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[38\]_B mprj_logic_high_inst/HI[368] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[76\] _538_/Y la_buf\[76\]/TE vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_29_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[24\]_A _422_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] user_to_mprj_in_gates\[65\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[65\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[29\]_B mprj_logic_high_inst/HI[359] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[5\]_A_N la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[1\]_A _591_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[99\]_TE la_buf\[99\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y vssd vssd vccd vccd la_data_in_mprj[35]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__501__A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[75\] la_iena_mprj[75] mprj_logic_high_inst/HI[405] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[75\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _362_/Y mprj_logic_high_inst/HI[303] vssd vssd vccd
+ vccd la_oenb_core[101] sky130_fd_sc_hd__einvp_8
X_600_ la_oenb_mprj[10] vssd vssd vccd vccd _600_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[31\] _621_/Y mprj_logic_high_inst/HI[233] vssd vssd vccd
+ vccd la_oenb_core[31] sky130_fd_sc_hd__einvp_8
X_531_ la_data_out_mprj[69] vssd vssd vccd vccd _531_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[53\] la_oenb_mprj[53] la_buf_enable\[53\]/B vssd vssd vccd vccd la_buf\[53\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[50\]_A_N la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_462_ la_data_out_mprj[0] vssd vssd vccd vccd _462_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_393_ mprj_we_o_core vssd vssd vccd vccd _393_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[39\] _501_/Y la_buf\[39\]/TE vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[65\]_A_N la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__411__A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[18\]_A_N la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] user_to_mprj_in_gates\[28\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[28\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[101\]_TE la_buf\[101\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[0\]_A _398_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[19\]_A _449_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[79\] _340_/Y mprj_logic_high_inst/HI[281] vssd vssd vccd
+ vccd la_oenb_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_2_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[27\] _457_/Y mprj_dat_buf\[27\]/TE vssd vssd vccd vccd mprj_dat_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[4\]_TE mprj_dat_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[0\]_B mprj_logic_high_inst/HI[330] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_514_ la_data_out_mprj[52] vssd vssd vccd vccd _514_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_445_ mprj_dat_o_core[15] vssd vssd vccd vccd _445_/Y sky130_fd_sc_hd__inv_2
X_376_ la_oenb_mprj[115] vssd vssd vccd vccd _376_/Y sky130_fd_sc_hd__inv_2
XANTENNA__406__A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[22\] _420_/Y mprj_adr_buf\[22\]/TE vssd vssd vccd vccd mprj_adr_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[121\]_B la_buf_enable\[121\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high_inst/HI[273] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[7\] la_oenb_mprj[7] la_buf_enable\[7\]/B vssd vssd vccd vccd la_buf\[7\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_9_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[112\]_B la_buf_enable\[112\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[38\] la_iena_mprj[38] mprj_logic_high_inst/HI[368] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[38\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[16\] la_oenb_mprj[16] la_buf_enable\[16\]/B vssd vssd vccd vccd la_buf\[16\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[121\] la_oenb_mprj[121] la_buf_enable\[121\]/B vssd vssd vccd vccd
+ la_buf\[121\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[6\]_A _468_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high_inst/HI[296] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[103\]_B la_buf_enable\[103\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_428_ mprj_adr_o_core[30] vssd vssd vccd vccd _428_/Y sky130_fd_sc_hd__inv_2
X_359_ la_oenb_mprj[98] vssd vssd vccd vccd _359_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] user_to_mprj_in_gates\[95\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[95\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[21\] _483_/Y la_buf\[21\]/TE vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__einvp_8
XFILLER_26_1403 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y vssd vssd vccd vccd la_data_in_mprj[65]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] user_to_mprj_in_gates\[10\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[10\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_30_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1863 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] user_to_mprj_in_gates\[121\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[121\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_2_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__504__A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[61\] _651_/Y mprj_logic_high_inst/HI[263] vssd vssd vccd
+ vccd la_oenb_core[61] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[83\] la_oenb_mprj[83] la_buf_enable\[83\]/B vssd vssd vccd vccd la_buf\[83\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[69\] _531_/Y la_buf\[69\]/TE vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__einvp_8
XFILLER_38_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__414__A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[125\] _587_/Y la_buf\[125\]/TE vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_26_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high_inst/HI[308] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] user_to_mprj_in_gates\[58\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[58\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_34_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[20\] la_iena_mprj[20] mprj_logic_high_inst/HI[350] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[20\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[106\]_A_N la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__409__A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y vssd vssd vccd vccd la_data_in_mprj[28]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[28\]_TE mprj_logic_high_inst/HI[230] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[0\]_B la_buf_enable\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[124\]_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[68\] la_iena_mprj[68] mprj_logic_high_inst/HI[398] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[68\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[115\]_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_530_ la_data_out_mprj[68] vssd vssd vccd vccd _530_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[6\] _596_/Y mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd la_oenb_core[6] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[24\] _614_/Y mprj_logic_high_inst/HI[226] vssd vssd vccd
+ vccd la_oenb_core[24] sky130_fd_sc_hd__einvp_8
X_461_ mprj_dat_o_core[31] vssd vssd vccd vccd _461_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[46\] la_oenb_mprj[46] la_buf_enable\[46\]/B vssd vssd vccd vccd la_buf\[46\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_13_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_392_ mprj_stb_o_core vssd vssd vccd vccd _392_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[4\]_A_N la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[106\]_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[15\]_TE mprj_dat_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__602__A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__512__A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[95\]_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_513_ la_data_out_mprj[51] vssd vssd vccd vccd _513_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_444_ mprj_dat_o_core[14] vssd vssd vccd vccd _444_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[51\] _513_/Y la_buf\[51\]/TE vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__einvp_8
X_375_ la_oenb_mprj[114] vssd vssd vccd vccd _375_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[123\] la_iena_mprj[123] mprj_logic_high_inst/HI[453] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[123\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__422__A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[15\] _413_/Y mprj_adr_buf\[15\]/TE vssd vssd vccd vccd mprj_adr_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y vssd vssd vccd vccd la_data_in_mprj[95]
+ sky130_fd_sc_hd__inv_8
XFILLER_27_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[86\]_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] user_to_mprj_in_gates\[40\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[40\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[10\]_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__332__A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] user_to_mprj_in_gates\[2\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[2\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[77\]_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[64\]_A_N la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[79\]_A_N la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__507__A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[91\] _352_/Y mprj_logic_high_inst/HI[293] vssd vssd vccd
+ vccd la_oenb_core[91] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[17\]_A_N la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[68\]_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[99\] _561_/Y la_buf\[99\]/TE vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[4\] la_iena_mprj[4] mprj_logic_high_inst/HI[334] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[4\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[114\] la_oenb_mprj[114] la_buf_enable\[114\]/B vssd vssd vccd vccd
+ la_buf\[114\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_1_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__417__A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_427_ mprj_adr_o_core[29] vssd vssd vccd vccd _427_/Y sky130_fd_sc_hd__inv_2
X_358_ la_oenb_mprj[97] vssd vssd vccd vccd _358_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y vssd vssd vccd vccd la_data_in_mprj[10]
+ sky130_fd_sc_hd__inv_8
XFILLER_6_794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] user_to_mprj_in_gates\[88\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[88\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[59\]_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_TE mprj_adr_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[50\] la_iena_mprj[50] mprj_logic_high_inst/HI[380] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[50\]/B sky130_fd_sc_hd__and2_1
XFILLER_9_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y vssd vssd vccd vccd la_data_in_mprj[2]
+ sky130_fd_sc_hd__inv_8
XFILLER_11_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[14\] _476_/Y la_buf\[14\]/TE vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_3_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[7\] _405_/Y mprj_adr_buf\[7\]/TE vssd vssd vccd vccd mprj_adr_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_18_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y vssd vssd vccd vccd la_data_in_mprj[58]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__610__A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] user_to_mprj_in_gates\[114\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[114\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[120\]_B user_to_mprj_in_gates\[120\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[98\] la_iena_mprj[98] mprj_logic_high_inst/HI[428] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[98\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high_inst/HI[286] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[124\] _385_/Y mprj_logic_high_inst/HI[326] vssd vssd vccd
+ vccd la_oenb_core[124] sky130_fd_sc_hd__einvp_8
XANTENNA__520__A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2160 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[54\] _644_/Y mprj_logic_high_inst/HI[256] vssd vssd vccd
+ vccd la_oenb_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_5_2254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[76\] la_oenb_mprj[76] la_buf_enable\[76\]/B vssd vssd vccd vccd la_buf\[76\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[118\] _580_/Y la_buf\[118\]/TE vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[111] sky130_fd_sc_hd__inv_8
XANTENNA__430__A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__605__A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__340__A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[13\] la_iena_mprj[13] mprj_logic_high_inst/HI[343] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[13\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[106\]_A _568_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__515__A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[81\] _543_/Y la_buf\[81\]/TE vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_1_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__425__A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[52\]_B la_buf_enable\[52\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] user_to_mprj_in_gates\[70\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[70\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[124\]_B mprj_logic_high_inst/HI[454] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_clk_buf _389_/Y mprj_clk_buf/TE vssd vssd vccd vccd user_clock sky130_fd_sc_hd__einvp_8
XFILLER_35_785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__335__A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[25\]_A _487_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[115\]_B mprj_logic_high_inst/HI[445] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_460_ mprj_dat_o_core[30] vssd vssd vccd vccd _460_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[17\] _607_/Y mprj_logic_high_inst/HI[219] vssd vssd vccd
+ vccd la_oenb_core[17] sky130_fd_sc_hd__einvp_8
X_391_ mprj_cyc_o_core vssd vssd vccd vccd _391_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[39\] la_oenb_mprj[39] la_buf_enable\[39\]/B vssd vssd vccd vccd la_buf\[39\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_13_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[16\]_A _478_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[34\]_B la_buf_enable\[34\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[3\]_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[106\]_B mprj_logic_high_inst/HI[436] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_589_ la_data_out_mprj[127] vssd vssd vccd vccd _589_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y vssd vssd vccd vccd la_data_in_mprj[40]
+ sky130_fd_sc_hd__inv_8
XFILLER_38_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[25\]_B la_buf_enable\[25\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[105\]_A_N la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high_inst/HI[321] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[16\]_B la_buf_enable\[16\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[80\] la_iena_mprj[80] mprj_logic_high_inst/HI[410] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[80\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_1196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[95\]_B mprj_logic_high_inst/HI[425] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_512_ la_data_out_mprj[50] vssd vssd vccd vccd _512_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_443_ mprj_dat_o_core[13] vssd vssd vccd vccd _443_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high_inst/HI[220] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[44\] _506_/Y la_buf\[44\]/TE vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__einvp_8
X_374_ la_oenb_mprj[113] vssd vssd vccd vccd _374_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[116\] la_iena_mprj[116] mprj_logic_high_inst/HI[446] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[116\]/B sky130_fd_sc_hd__and2_1
XFILLER_9_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[100\] _562_/Y la_buf\[100\]/TE vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[86\]_B mprj_logic_high_inst/HI[416] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y vssd vssd vccd vccd la_data_in_mprj[88]
+ sky130_fd_sc_hd__inv_8
XFILLER_24_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] user_to_mprj_in_gates\[33\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[33\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[10\]_B mprj_logic_high_inst/HI[340] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__613__A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[3\]_A_N la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__523__A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[84\] _345_/Y mprj_logic_high_inst/HI[286] vssd vssd vccd
+ vccd la_oenb_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[107\] la_oenb_mprj[107] la_buf_enable\[107\]/B vssd vssd vccd vccd
+ la_buf\[107\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_2_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_426_ mprj_adr_o_core[28] vssd vssd vccd vccd _426_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_357_ la_oenb_mprj[96] vssd vssd vccd vccd _357_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__433__A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[59\]_B mprj_logic_high_inst/HI[389] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__608__A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__343__A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[43\] la_iena_mprj[43] mprj_logic_high_inst/HI[373] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[43\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__518__A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[7\]_TE mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[21\] la_oenb_mprj[21] la_buf_enable\[21\]/B vssd vssd vccd vccd la_buf\[21\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__428__A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_409_ mprj_adr_o_core[11] vssd vssd vccd vccd _409_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_1409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[63\]_A_N la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[27\]_A _425_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[78\]_A_N la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_sel_buf\[2\]_TE mprj_sel_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] user_to_mprj_in_gates\[107\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[107\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__338__A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[16\]_A_N la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[4\]_A _594_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[18\]_A _416_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[117\] _378_/Y mprj_logic_high_inst/HI[319] vssd vssd vccd
+ vccd la_oenb_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_7_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_931 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[47\] _637_/Y mprj_logic_high_inst/HI[249] vssd vssd vccd
+ vccd la_oenb_core[47] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[69\] la_oenb_mprj[69] la_buf_enable\[69\]/B vssd vssd vccd vccd la_buf\[69\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[104] sky130_fd_sc_hd__inv_8
XFILLER_38_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y vssd vssd vccd vccd la_data_in_mprj[70]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[104\]_TE la_buf\[104\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__621__A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[3\] _433_/Y mprj_dat_buf\[3\]/TE vssd vssd vccd vccd mprj_dat_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_38_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__531__A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[74\] _536_/Y la_buf\[74\]/TE vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__einvp_8
XFILLER_1_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__441__A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] user_to_mprj_in_gates\[63\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[63\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high_inst/HI[276] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__616__A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[3\]_A _401_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__351__A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_390_ caravel_clk2 vssd vssd vccd vccd _390_/Y sky130_fd_sc_hd__inv_2
XANTENNA__526__A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[3\]_B mprj_logic_high_inst/HI[333] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high_inst/HI[299] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_657_ la_oenb_mprj[67] vssd vssd vccd vccd _657_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_588_ la_data_out_mprj[126] vssd vssd vccd vccd _588_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__436__A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y vssd vssd vccd vccd la_data_in_mprj[33]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[124\]_B la_buf_enable\[124\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__346__A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[73\] la_iena_mprj[73] mprj_logic_high_inst/HI[403] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[73\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[115\]_B la_buf_enable\[115\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_511_ la_data_out_mprj[49] vssd vssd vccd vccd _511_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[51\] la_oenb_mprj[51] la_buf_enable\[51\]/B vssd vssd vccd vccd la_buf\[51\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_442_ mprj_dat_o_core[12] vssd vssd vccd vccd _442_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_373_ la_oenb_mprj[112] vssd vssd vccd vccd _373_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[37\] _499_/Y la_buf\[37\]/TE vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__einvp_8
XFILLER_35_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[109\] la_iena_mprj[109] mprj_logic_high_inst/HI[439] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[109\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[9\]_A _471_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[106\]_B la_buf_enable\[106\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] user_to_mprj_in_gates\[26\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[26\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[77\] _338_/Y mprj_logic_high_inst/HI[279] vssd vssd vccd
+ vccd la_oenb_core[77] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[99\] la_oenb_mprj[99] la_buf_enable\[99\]/B vssd vssd vccd vccd la_buf\[99\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[25\] _455_/Y mprj_dat_buf\[25\]/TE vssd vssd vccd vccd mprj_dat_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_425_ mprj_adr_o_core[27] vssd vssd vccd vccd _425_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[104\]_A_N la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_356_ la_oenb_mprj[95] vssd vssd vccd vccd _356_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[20\] _418_/Y mprj_adr_buf\[20\]/TE vssd vssd vccd vccd mprj_adr_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[119\]_A_N la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high_inst/HI[311] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__624__A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[5\] la_oenb_mprj[5] la_buf_enable\[5\]/B vssd vssd vccd vccd la_buf\[5\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_TE la_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[36\] la_iena_mprj[36] mprj_logic_high_inst/HI[366] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[36\]/B sky130_fd_sc_hd__and2_1
XFILLER_23_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__534__A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[14\] la_oenb_mprj[14] la_buf_enable\[14\]/B vssd vssd vccd vccd la_buf\[14\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_7_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_408_ mprj_adr_o_core[10] vssd vssd vccd vccd _408_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__444__A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_339_ la_oenb_mprj[78] vssd vssd vccd vccd _339_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] user_to_mprj_in_gates\[93\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[93\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[2\]_A_N la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1826 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__619__A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__354__A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__529__A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__439__A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y vssd vssd vccd vccd la_data_in_mprj[63]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[18\]_TE mprj_dat_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[3\]_B la_buf_enable\[3\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[127\]_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__349__A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[81\] la_oenb_mprj[81] la_buf_enable\[81\]/B vssd vssd vccd vccd la_buf\[81\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[118\]_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[62\]_A_N la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[67\] _529_/Y la_buf\[67\]/TE vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__einvp_8
XFILLER_16_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[77\]_A_N la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[123\] _585_/Y la_buf\[123\]/TE vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[15\]_A_N la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[109\]_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] user_to_mprj_in_gates\[56\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[56\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[40\]_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__632__A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__542__A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[98\]_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_656_ la_oenb_mprj[66] vssd vssd vccd vccd _656_/Y sky130_fd_sc_hd__inv_2
X_587_ la_data_out_mprj[125] vssd vssd vccd vccd _587_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[22\]_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y vssd vssd vccd vccd la_data_in_mprj[26]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__452__A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[89\]_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[41\]_TE mprj_logic_high_inst/HI[243] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__627__A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[13\]_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__362__A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[66\] la_iena_mprj[66] mprj_logic_high_inst/HI[396] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[66\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_510_ la_data_out_mprj[48] vssd vssd vccd vccd _510_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[0\]_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__537__A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[22\] _612_/Y mprj_logic_high_inst/HI[224] vssd vssd vccd
+ vccd la_oenb_core[22] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[4\] _594_/Y mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd la_oenb_core[4] sky130_fd_sc_hd__einvp_8
X_441_ mprj_dat_o_core[11] vssd vssd vccd vccd _441_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[44\] la_oenb_mprj[44] la_buf_enable\[44\]/B vssd vssd vccd vccd la_buf\[44\]/TE
+ sky130_fd_sc_hd__and2b_1
X_372_ la_oenb_mprj[111] vssd vssd vccd vccd _372_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[64\]_TE mprj_logic_high_inst/HI[266] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__447__A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_639_ la_oenb_mprj[49] vssd vssd vccd vccd _639_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] user_to_mprj_in_gates\[19\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[19\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__357__A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high_inst/HI[289] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1586 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[18\] _448_/Y mprj_dat_buf\[18\]/TE vssd vssd vccd vccd mprj_dat_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XFILLER_18_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_424_ mprj_adr_o_core[26] vssd vssd vccd vccd _424_/Y sky130_fd_sc_hd__inv_2
X_355_ la_oenb_mprj[94] vssd vssd vccd vccd _355_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[121\] la_iena_mprj[121] mprj_logic_high_inst/HI[451] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[121\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[13\] _411_/Y mprj_adr_buf\[13\]/TE vssd vssd vccd vccd mprj_adr_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[127] sky130_fd_sc_hd__inv_8
XFILLER_29_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y vssd vssd vccd vccd la_data_in_mprj[93]
+ sky130_fd_sc_hd__inv_8
XFILLER_36_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[82\]_A _544_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__640__A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] user_to_mprj_in_gates\[0\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[0\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[29\] la_iena_mprj[29] mprj_logic_high_inst/HI[359] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[29\]/B sky130_fd_sc_hd__and2_1
XFILLER_23_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[123\]_B user_to_mprj_in_gates\[123\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[91\]_B la_buf_enable\[91\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__550__A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[97\] _559_/Y la_buf\[97\]/TE vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[2\] la_iena_mprj[2] mprj_logic_high_inst/HI[332] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[2\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[112\] la_oenb_mprj[112] la_buf_enable\[112\]/B vssd vssd vccd vccd
+ la_buf\[112\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[127\]_A _589_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_407_ mprj_adr_o_core[9] vssd vssd vccd vccd _407_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[114\]_B user_to_mprj_in_gates\[114\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_338_ la_oenb_mprj[77] vssd vssd vccd vccd _338_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[64\]_A _526_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[82\]_B la_buf_enable\[82\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__460__A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] user_to_mprj_in_gates\[86\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[86\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__635__A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__370__A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[103\]_A_N la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[118\]_A_N la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y vssd vssd vccd vccd la_data_in_mprj[0]
+ sky130_fd_sc_hd__inv_8
XANTENNA__545__A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[64\]_B la_buf_enable\[64\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[8\] _470_/Y la_buf\[8\]/TE vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__einvp_8
Xla_buf\[12\] _474_/Y la_buf\[12\]/TE vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__einvp_8
XFILLER_3_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[5\] _403_/Y mprj_adr_buf\[5\]/TE vssd vssd vccd vccd mprj_adr_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_35_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y vssd vssd vccd vccd la_data_in_mprj[56]
+ sky130_fd_sc_hd__inv_8
XANTENNA__455__A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[55\]_B la_buf_enable\[55\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[127\]_B mprj_logic_high_inst/HI[457] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_2336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] user_to_mprj_in_gates\[112\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[112\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__365__A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[46\]_B la_buf_enable\[46\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[96\] la_iena_mprj[96] mprj_logic_high_inst/HI[426] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[96\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[122\] _383_/Y mprj_logic_high_inst/HI[324] vssd vssd vccd
+ vccd la_oenb_core[122] sky130_fd_sc_hd__einvp_8
XFILLER_27_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[3\] _397_/Y mprj_sel_buf\[3\]/TE vssd vssd vccd vccd mprj_sel_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[118\]_B mprj_logic_high_inst/HI[448] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[52\] _642_/Y mprj_logic_high_inst/HI[254] vssd vssd vccd
+ vccd la_oenb_core[52] sky130_fd_sc_hd__einvp_8
XFILLER_5_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[74\] la_oenb_mprj[74] la_buf_enable\[74\]/B vssd vssd vccd vccd la_buf\[74\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[1\]_A_N la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[19\]_A _481_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[37\]_B la_buf_enable\[37\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[6\]_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[116\] _578_/Y la_buf\[116\]/TE vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_3_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_clk2_buf_A _390_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[109\]_B mprj_logic_high_inst/HI[439] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] user_to_mprj_in_gates\[49\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[49\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[40\]_B mprj_logic_high_inst/HI[370] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_B la_buf_enable\[28\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[11\] la_iena_mprj[11] mprj_logic_high_inst/HI[341] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[11\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_B mprj_logic_high_inst/HI[361] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[19\]_B la_buf_enable\[19\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[98\]_B mprj_logic_high_inst/HI[428] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_655_ la_oenb_mprj[65] vssd vssd vccd vccd _655_/Y sky130_fd_sc_hd__inv_2
X_586_ la_data_out_mprj[124] vssd vssd vccd vccd _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[22\]_B mprj_logic_high_inst/HI[352] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y vssd vssd vccd vccd la_data_in_mprj[19]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_oen_buffers\[12\]_A _602_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[89\]_B mprj_logic_high_inst/HI[419] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[13\]_B mprj_logic_high_inst/HI[343] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__643__A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[61\]_A_N la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[76\]_A_N la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[59\] la_iena_mprj[59] mprj_logic_high_inst/HI[389] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[59\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_2182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_irq_ena_buf\[0\]_B user_irq_ena_buf\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_440_ mprj_dat_o_core[10] vssd vssd vccd vccd _440_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[15\] _605_/Y mprj_logic_high_inst/HI[217] vssd vssd vccd
+ vccd la_oenb_core[15] sky130_fd_sc_hd__einvp_8
X_371_ la_oenb_mprj[110] vssd vssd vccd vccd _371_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[37\] la_oenb_mprj[37] la_buf_enable\[37\]/B vssd vssd vccd vccd la_buf\[37\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[14\]_A_N la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__553__A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[29\]_A_N la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_638_ la_oenb_mprj[48] vssd vssd vccd vccd _638_/Y sky130_fd_sc_hd__inv_2
X_569_ la_data_out_mprj[107] vssd vssd vccd vccd _569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__463__A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__638__A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__373__A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__548__A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_423_ mprj_adr_o_core[25] vssd vssd vccd vccd _423_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_A _451_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[42\] _504_/Y la_buf\[42\]/TE vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__einvp_8
X_354_ la_oenb_mprj[93] vssd vssd vccd vccd _354_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[114\] la_iena_mprj[114] mprj_logic_high_inst/HI[444] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[114\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y vssd vssd vccd vccd la_data_in_mprj[86]
+ sky130_fd_sc_hd__inv_8
XFILLER_36_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__458__A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[107\]_TE la_buf\[107\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] user_to_mprj_in_gates\[31\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[31\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[12\]_A _442_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[6\]_TE mprj_adr_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__368__A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[82\] _343_/Y mprj_logic_high_inst/HI[284] vssd vssd vccd
+ vccd la_oenb_core[82] sky130_fd_sc_hd__einvp_8
XFILLER_10_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[30\] _460_/Y mprj_dat_buf\[30\]/TE vssd vssd vccd vccd mprj_dat_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[105\] la_oenb_mprj[105] la_buf_enable\[105\]/B vssd vssd vccd vccd
+ la_buf\[105\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_18_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_406_ mprj_adr_o_core[8] vssd vssd vccd vccd _406_/Y sky130_fd_sc_hd__inv_2
X_337_ la_oenb_mprj[76] vssd vssd vccd vccd _337_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] user_to_mprj_in_gates\[79\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[79\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high_inst/HI[279] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__651__A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[41\] la_iena_mprj[41] mprj_logic_high_inst/HI[371] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[41\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__561__A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1710 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y vssd vssd vccd vccd la_data_in_mprj[49]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__471__A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] user_to_mprj_in_gates\[105\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[105\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__646__A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_logic_high_inst mprj2_pwrgood/A vccd2 vssd mprj2_logic_high
XANTENNA_mprj_adr_buf\[6\]_A _404_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__381__A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[89\] la_iena_mprj[89] mprj_logic_high_inst/HI[419] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[89\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[115\] _376_/Y mprj_logic_high_inst/HI[317] vssd vssd vccd
+ vccd la_oenb_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_5_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[45\] _635_/Y mprj_logic_high_inst/HI[247] vssd vssd vccd
+ vccd la_oenb_core[45] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[67\] la_oenb_mprj[67] la_buf_enable\[67\]/B vssd vssd vccd vccd la_buf\[67\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__556__A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[6\]_B mprj_logic_high_inst/HI[336] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[109\] _571_/Y la_buf\[109\]/TE vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_3_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[102] sky130_fd_sc_hd__inv_8
XFILLER_6_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__466__A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[102\]_A_N la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[117\]_A_N la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[127\]_B la_buf_enable\[127\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[1\] _431_/Y mprj_dat_buf\[1\]/TE vssd vssd vccd vccd mprj_dat_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_logic_high_inst mprj_rstn_buf/TE la_buf_enable\[26\]/B la_buf_enable\[27\]/B
+ la_buf_enable\[28\]/B la_buf_enable\[29\]/B la_buf_enable\[30\]/B la_buf_enable\[31\]/B
+ la_buf_enable\[32\]/B la_buf_enable\[33\]/B la_buf_enable\[34\]/B la_buf_enable\[35\]/B
+ mprj_adr_buf\[0\]/TE la_buf_enable\[36\]/B la_buf_enable\[37\]/B la_buf_enable\[38\]/B
+ la_buf_enable\[39\]/B la_buf_enable\[40\]/B la_buf_enable\[41\]/B la_buf_enable\[42\]/B
+ la_buf_enable\[43\]/B la_buf_enable\[44\]/B la_buf_enable\[45\]/B mprj_adr_buf\[1\]/TE
+ la_buf_enable\[46\]/B la_buf_enable\[47\]/B la_buf_enable\[48\]/B la_buf_enable\[49\]/B
+ la_buf_enable\[50\]/B la_buf_enable\[51\]/B la_buf_enable\[52\]/B la_buf_enable\[53\]/B
+ la_buf_enable\[54\]/B la_buf_enable\[55\]/B mprj_adr_buf\[2\]/TE la_buf_enable\[56\]/B
+ la_buf_enable\[57\]/B la_buf_enable\[58\]/B la_buf_enable\[59\]/B la_buf_enable\[60\]/B
+ la_buf_enable\[61\]/B la_buf_enable\[62\]/B la_buf_enable\[63\]/B la_buf_enable\[64\]/B
+ la_buf_enable\[65\]/B mprj_adr_buf\[3\]/TE la_buf_enable\[66\]/B la_buf_enable\[67\]/B
+ la_buf_enable\[68\]/B la_buf_enable\[69\]/B la_buf_enable\[70\]/B la_buf_enable\[71\]/B
+ la_buf_enable\[72\]/B la_buf_enable\[73\]/B la_buf_enable\[74\]/B la_buf_enable\[75\]/B
+ mprj_adr_buf\[4\]/TE la_buf_enable\[76\]/B la_buf_enable\[77\]/B la_buf_enable\[78\]/B
+ la_buf_enable\[79\]/B la_buf_enable\[80\]/B la_buf_enable\[81\]/B la_buf_enable\[82\]/B
+ la_buf_enable\[83\]/B la_buf_enable\[84\]/B la_buf_enable\[85\]/B mprj_adr_buf\[5\]/TE
+ la_buf_enable\[86\]/B la_buf_enable\[87\]/B la_buf_enable\[88\]/B la_buf_enable\[89\]/B
+ la_buf_enable\[90\]/B la_buf_enable\[91\]/B la_buf_enable\[92\]/B la_buf_enable\[93\]/B
+ la_buf_enable\[94\]/B la_buf_enable\[95\]/B mprj_adr_buf\[6\]/TE la_buf_enable\[96\]/B
+ la_buf_enable\[97\]/B la_buf_enable\[98\]/B la_buf_enable\[99\]/B la_buf_enable\[100\]/B
+ la_buf_enable\[101\]/B la_buf_enable\[102\]/B la_buf_enable\[103\]/B la_buf_enable\[104\]/B
+ la_buf_enable\[105\]/B mprj_adr_buf\[7\]/TE la_buf_enable\[106\]/B la_buf_enable\[107\]/B
+ la_buf_enable\[108\]/B la_buf_enable\[109\]/B la_buf_enable\[110\]/B la_buf_enable\[111\]/B
+ la_buf_enable\[112\]/B la_buf_enable\[113\]/B la_buf_enable\[114\]/B la_buf_enable\[115\]/B
+ mprj_adr_buf\[8\]/TE la_buf_enable\[116\]/B la_buf_enable\[117\]/B la_buf_enable\[118\]/B
+ la_buf_enable\[119\]/B la_buf_enable\[120\]/B la_buf_enable\[121\]/B la_buf_enable\[122\]/B
+ la_buf_enable\[123\]/B la_buf_enable\[124\]/B mprj_adr_buf\[9\]/TE mprj_clk_buf/TE
+ la_buf_enable\[126\]/B la_buf_enable\[127\]/B mprj_logic_high_inst/HI[202] mprj_logic_high_inst/HI[203]
+ mprj_logic_high_inst/HI[204] mprj_logic_high_inst/HI[205] mprj_logic_high_inst/HI[206]
+ mprj_logic_high_inst/HI[207] mprj_logic_high_inst/HI[208] mprj_logic_high_inst/HI[209]
+ mprj_adr_buf\[10\]/TE mprj_logic_high_inst/HI[210] mprj_logic_high_inst/HI[211]
+ mprj_logic_high_inst/HI[212] mprj_logic_high_inst/HI[213] mprj_logic_high_inst/HI[214]
+ mprj_logic_high_inst/HI[215] mprj_logic_high_inst/HI[216] mprj_logic_high_inst/HI[217]
+ mprj_logic_high_inst/HI[218] mprj_logic_high_inst/HI[219] mprj_adr_buf\[11\]/TE
+ mprj_logic_high_inst/HI[220] mprj_logic_high_inst/HI[221] mprj_logic_high_inst/HI[222]
+ mprj_logic_high_inst/HI[223] mprj_logic_high_inst/HI[224] mprj_logic_high_inst/HI[225]
+ mprj_logic_high_inst/HI[226] mprj_logic_high_inst/HI[227] mprj_logic_high_inst/HI[228]
+ mprj_logic_high_inst/HI[229] mprj_adr_buf\[12\]/TE mprj_logic_high_inst/HI[230]
+ mprj_logic_high_inst/HI[231] mprj_logic_high_inst/HI[232] mprj_logic_high_inst/HI[233]
+ mprj_logic_high_inst/HI[234] mprj_logic_high_inst/HI[235] mprj_logic_high_inst/HI[236]
+ mprj_logic_high_inst/HI[237] mprj_logic_high_inst/HI[238] mprj_logic_high_inst/HI[239]
+ mprj_adr_buf\[13\]/TE mprj_logic_high_inst/HI[240] mprj_logic_high_inst/HI[241]
+ mprj_logic_high_inst/HI[242] mprj_logic_high_inst/HI[243] mprj_logic_high_inst/HI[244]
+ mprj_logic_high_inst/HI[245] mprj_logic_high_inst/HI[246] mprj_logic_high_inst/HI[247]
+ mprj_logic_high_inst/HI[248] mprj_logic_high_inst/HI[249] mprj_adr_buf\[14\]/TE
+ mprj_logic_high_inst/HI[250] mprj_logic_high_inst/HI[251] mprj_logic_high_inst/HI[252]
+ mprj_logic_high_inst/HI[253] mprj_logic_high_inst/HI[254] mprj_logic_high_inst/HI[255]
+ mprj_logic_high_inst/HI[256] mprj_logic_high_inst/HI[257] mprj_logic_high_inst/HI[258]
+ mprj_logic_high_inst/HI[259] mprj_adr_buf\[15\]/TE mprj_logic_high_inst/HI[260]
+ mprj_logic_high_inst/HI[261] mprj_logic_high_inst/HI[262] mprj_logic_high_inst/HI[263]
+ mprj_logic_high_inst/HI[264] mprj_logic_high_inst/HI[265] mprj_logic_high_inst/HI[266]
+ mprj_logic_high_inst/HI[267] mprj_logic_high_inst/HI[268] mprj_logic_high_inst/HI[269]
+ mprj_adr_buf\[16\]/TE mprj_logic_high_inst/HI[270] mprj_logic_high_inst/HI[271]
+ mprj_logic_high_inst/HI[272] mprj_logic_high_inst/HI[273] mprj_logic_high_inst/HI[274]
+ mprj_logic_high_inst/HI[275] mprj_logic_high_inst/HI[276] mprj_logic_high_inst/HI[277]
+ mprj_logic_high_inst/HI[278] mprj_logic_high_inst/HI[279] mprj_adr_buf\[17\]/TE
+ mprj_logic_high_inst/HI[280] mprj_logic_high_inst/HI[281] mprj_logic_high_inst/HI[282]
+ mprj_logic_high_inst/HI[283] mprj_logic_high_inst/HI[284] mprj_logic_high_inst/HI[285]
+ mprj_logic_high_inst/HI[286] mprj_logic_high_inst/HI[287] mprj_logic_high_inst/HI[288]
+ mprj_logic_high_inst/HI[289] mprj_adr_buf\[18\]/TE mprj_logic_high_inst/HI[290]
+ mprj_logic_high_inst/HI[291] mprj_logic_high_inst/HI[292] mprj_logic_high_inst/HI[293]
+ mprj_logic_high_inst/HI[294] mprj_logic_high_inst/HI[295] mprj_logic_high_inst/HI[296]
+ mprj_logic_high_inst/HI[297] mprj_logic_high_inst/HI[298] mprj_logic_high_inst/HI[299]
+ mprj_adr_buf\[19\]/TE mprj_clk2_buf/TE mprj_logic_high_inst/HI[300] mprj_logic_high_inst/HI[301]
+ mprj_logic_high_inst/HI[302] mprj_logic_high_inst/HI[303] mprj_logic_high_inst/HI[304]
+ mprj_logic_high_inst/HI[305] mprj_logic_high_inst/HI[306] mprj_logic_high_inst/HI[307]
+ mprj_logic_high_inst/HI[308] mprj_logic_high_inst/HI[309] mprj_adr_buf\[20\]/TE
+ mprj_logic_high_inst/HI[310] mprj_logic_high_inst/HI[311] mprj_logic_high_inst/HI[312]
+ mprj_logic_high_inst/HI[313] mprj_logic_high_inst/HI[314] mprj_logic_high_inst/HI[315]
+ mprj_logic_high_inst/HI[316] mprj_logic_high_inst/HI[317] mprj_logic_high_inst/HI[318]
+ mprj_logic_high_inst/HI[319] mprj_adr_buf\[21\]/TE mprj_logic_high_inst/HI[320]
+ mprj_logic_high_inst/HI[321] mprj_logic_high_inst/HI[322] mprj_logic_high_inst/HI[323]
+ mprj_logic_high_inst/HI[324] mprj_logic_high_inst/HI[325] mprj_logic_high_inst/HI[326]
+ mprj_logic_high_inst/HI[327] mprj_logic_high_inst/HI[328] mprj_logic_high_inst/HI[329]
+ mprj_adr_buf\[22\]/TE mprj_logic_high_inst/HI[330] mprj_logic_high_inst/HI[331]
+ mprj_logic_high_inst/HI[332] mprj_logic_high_inst/HI[333] mprj_logic_high_inst/HI[334]
+ mprj_logic_high_inst/HI[335] mprj_logic_high_inst/HI[336] mprj_logic_high_inst/HI[337]
+ mprj_logic_high_inst/HI[338] mprj_logic_high_inst/HI[339] mprj_adr_buf\[23\]/TE
+ mprj_logic_high_inst/HI[340] mprj_logic_high_inst/HI[341] mprj_logic_high_inst/HI[342]
+ mprj_logic_high_inst/HI[343] mprj_logic_high_inst/HI[344] mprj_logic_high_inst/HI[345]
+ mprj_logic_high_inst/HI[346] mprj_logic_high_inst/HI[347] mprj_logic_high_inst/HI[348]
+ mprj_logic_high_inst/HI[349] mprj_adr_buf\[24\]/TE mprj_logic_high_inst/HI[350]
+ mprj_logic_high_inst/HI[351] mprj_logic_high_inst/HI[352] mprj_logic_high_inst/HI[353]
+ mprj_logic_high_inst/HI[354] mprj_logic_high_inst/HI[355] mprj_logic_high_inst/HI[356]
+ mprj_logic_high_inst/HI[357] mprj_logic_high_inst/HI[358] mprj_logic_high_inst/HI[359]
+ mprj_adr_buf\[25\]/TE mprj_logic_high_inst/HI[360] mprj_logic_high_inst/HI[361]
+ mprj_logic_high_inst/HI[362] mprj_logic_high_inst/HI[363] mprj_logic_high_inst/HI[364]
+ mprj_logic_high_inst/HI[365] mprj_logic_high_inst/HI[366] mprj_logic_high_inst/HI[367]
+ mprj_logic_high_inst/HI[368] mprj_logic_high_inst/HI[369] mprj_adr_buf\[26\]/TE
+ mprj_logic_high_inst/HI[370] mprj_logic_high_inst/HI[371] mprj_logic_high_inst/HI[372]
+ mprj_logic_high_inst/HI[373] mprj_logic_high_inst/HI[374] mprj_logic_high_inst/HI[375]
+ mprj_logic_high_inst/HI[376] mprj_logic_high_inst/HI[377] mprj_logic_high_inst/HI[378]
+ mprj_logic_high_inst/HI[379] mprj_adr_buf\[27\]/TE mprj_logic_high_inst/HI[380]
+ mprj_logic_high_inst/HI[381] mprj_logic_high_inst/HI[382] mprj_logic_high_inst/HI[383]
+ mprj_logic_high_inst/HI[384] mprj_logic_high_inst/HI[385] mprj_logic_high_inst/HI[386]
+ mprj_logic_high_inst/HI[387] mprj_logic_high_inst/HI[388] mprj_logic_high_inst/HI[389]
+ mprj_adr_buf\[28\]/TE mprj_logic_high_inst/HI[390] mprj_logic_high_inst/HI[391]
+ mprj_logic_high_inst/HI[392] mprj_logic_high_inst/HI[393] mprj_logic_high_inst/HI[394]
+ mprj_logic_high_inst/HI[395] mprj_logic_high_inst/HI[396] mprj_logic_high_inst/HI[397]
+ mprj_logic_high_inst/HI[398] mprj_logic_high_inst/HI[399] mprj_adr_buf\[29\]/TE
+ mprj_cyc_buf/TE mprj_logic_high_inst/HI[400] mprj_logic_high_inst/HI[401] mprj_logic_high_inst/HI[402]
+ mprj_logic_high_inst/HI[403] mprj_logic_high_inst/HI[404] mprj_logic_high_inst/HI[405]
+ mprj_logic_high_inst/HI[406] mprj_logic_high_inst/HI[407] mprj_logic_high_inst/HI[408]
+ mprj_logic_high_inst/HI[409] mprj_adr_buf\[30\]/TE mprj_logic_high_inst/HI[410]
+ mprj_logic_high_inst/HI[411] mprj_logic_high_inst/HI[412] mprj_logic_high_inst/HI[413]
+ mprj_logic_high_inst/HI[414] mprj_logic_high_inst/HI[415] mprj_logic_high_inst/HI[416]
+ mprj_logic_high_inst/HI[417] mprj_logic_high_inst/HI[418] mprj_logic_high_inst/HI[419]
+ mprj_adr_buf\[31\]/TE mprj_logic_high_inst/HI[420] mprj_logic_high_inst/HI[421]
+ mprj_logic_high_inst/HI[422] mprj_logic_high_inst/HI[423] mprj_logic_high_inst/HI[424]
+ mprj_logic_high_inst/HI[425] mprj_logic_high_inst/HI[426] mprj_logic_high_inst/HI[427]
+ mprj_logic_high_inst/HI[428] mprj_logic_high_inst/HI[429] mprj_dat_buf\[0\]/TE mprj_logic_high_inst/HI[430]
+ mprj_logic_high_inst/HI[431] mprj_logic_high_inst/HI[432] mprj_logic_high_inst/HI[433]
+ mprj_logic_high_inst/HI[434] mprj_logic_high_inst/HI[435] mprj_logic_high_inst/HI[436]
+ mprj_logic_high_inst/HI[437] mprj_logic_high_inst/HI[438] mprj_logic_high_inst/HI[439]
+ mprj_dat_buf\[1\]/TE mprj_logic_high_inst/HI[440] mprj_logic_high_inst/HI[441] mprj_logic_high_inst/HI[442]
+ mprj_logic_high_inst/HI[443] mprj_logic_high_inst/HI[444] mprj_logic_high_inst/HI[445]
+ mprj_logic_high_inst/HI[446] mprj_logic_high_inst/HI[447] mprj_logic_high_inst/HI[448]
+ mprj_logic_high_inst/HI[449] mprj_dat_buf\[2\]/TE mprj_logic_high_inst/HI[450] mprj_logic_high_inst/HI[451]
+ mprj_logic_high_inst/HI[452] mprj_logic_high_inst/HI[453] mprj_logic_high_inst/HI[454]
+ mprj_logic_high_inst/HI[455] mprj_logic_high_inst/HI[456] mprj_logic_high_inst/HI[457]
+ user_irq_ena_buf\[0\]/B user_irq_ena_buf\[1\]/B mprj_dat_buf\[3\]/TE user_irq_ena_buf\[2\]/B
+ mprj_pwrgood/A mprj_dat_buf\[4\]/TE mprj_dat_buf\[5\]/TE mprj_dat_buf\[6\]/TE mprj_dat_buf\[7\]/TE
+ mprj_stb_buf/TE mprj_dat_buf\[8\]/TE mprj_dat_buf\[9\]/TE mprj_dat_buf\[10\]/TE
+ mprj_dat_buf\[11\]/TE mprj_dat_buf\[12\]/TE mprj_dat_buf\[13\]/TE mprj_dat_buf\[14\]/TE
+ mprj_dat_buf\[15\]/TE mprj_dat_buf\[16\]/TE mprj_dat_buf\[17\]/TE mprj_we_buf/TE
+ mprj_dat_buf\[18\]/TE mprj_dat_buf\[19\]/TE mprj_dat_buf\[20\]/TE mprj_dat_buf\[21\]/TE
+ mprj_dat_buf\[22\]/TE mprj_dat_buf\[23\]/TE mprj_dat_buf\[24\]/TE mprj_dat_buf\[25\]/TE
+ mprj_dat_buf\[26\]/TE mprj_dat_buf\[27\]/TE mprj_sel_buf\[0\]/TE mprj_dat_buf\[28\]/TE
+ mprj_dat_buf\[29\]/TE mprj_dat_buf\[30\]/TE mprj_dat_buf\[31\]/TE la_buf_enable\[0\]/B
+ la_buf_enable\[1\]/B la_buf_enable\[2\]/B la_buf_enable\[3\]/B la_buf_enable\[4\]/B
+ la_buf_enable\[5\]/B mprj_sel_buf\[1\]/TE la_buf_enable\[6\]/B la_buf_enable\[7\]/B
+ la_buf_enable\[8\]/B la_buf_enable\[9\]/B la_buf_enable\[10\]/B la_buf_enable\[11\]/B
+ la_buf_enable\[12\]/B la_buf_enable\[13\]/B la_buf_enable\[14\]/B la_buf_enable\[15\]/B
+ mprj_sel_buf\[2\]/TE la_buf_enable\[16\]/B la_buf_enable\[17\]/B la_buf_enable\[18\]/B
+ la_buf_enable\[19\]/B la_buf_enable\[20\]/B la_buf_enable\[21\]/B la_buf_enable\[22\]/B
+ la_buf_enable\[23\]/B la_buf_enable\[24\]/B la_buf_enable\[25\]/B mprj_sel_buf\[3\]/TE
+ vccd1 vssd la_buf_enable\[125\]/B mprj_logic_high
XFILLER_26_2292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__376__A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[118\]_B la_buf_enable\[118\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_654_ la_oenb_mprj[64] vssd vssd vccd vccd _654_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[72\] _534_/Y la_buf\[72\]/TE vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__einvp_8
XFILLER_29_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_585_ la_data_out_mprj[123] vssd vssd vccd vccd _585_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[109\]_B la_buf_enable\[109\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] user_to_mprj_in_gates\[61\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[61\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_TE la_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[0\]_A_N la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_370_ la_oenb_mprj[109] vssd vssd vccd vccd _370_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1439 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_637_ la_oenb_mprj[47] vssd vssd vccd vccd _637_/Y sky130_fd_sc_hd__inv_2
X_568_ la_data_out_mprj[106] vssd vssd vccd vccd _568_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y vssd vssd vccd vccd la_data_in_mprj[31]
+ sky130_fd_sc_hd__inv_8
X_499_ la_data_out_mprj[37] vssd vssd vccd vccd _499_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__654__A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[71\] la_iena_mprj[71] mprj_logic_high_inst/HI[401] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[71\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_422_ mprj_adr_o_core[24] vssd vssd vccd vccd _422_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__564__A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_353_ la_oenb_mprj[92] vssd vssd vccd vccd _353_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[35\] _497_/Y la_buf\[35\]/TE vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__einvp_8
XFILLER_35_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[107\] la_iena_mprj[107] mprj_logic_high_inst/HI[437] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[107\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y vssd vssd vccd vccd la_data_in_mprj[79]
+ sky130_fd_sc_hd__inv_8
XFILLER_24_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[60\]_A_N la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__474__A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] user_to_mprj_in_gates\[24\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[24\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[75\]_A_N la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[13\]_A_N la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__649__A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_A_N la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__384__A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[75\] _336_/Y mprj_logic_high_inst/HI[277] vssd vssd vccd
+ vccd la_oenb_core[75] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[97\] la_oenb_mprj[97] la_buf_enable\[97\]/B vssd vssd vccd vccd la_buf\[97\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[23\] _453_/Y mprj_dat_buf\[23\]/TE vssd vssd vccd vccd mprj_dat_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__559__A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_405_ mprj_adr_o_core[7] vssd vssd vccd vccd _405_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_336_ la_oenb_mprj[75] vssd vssd vccd vccd _336_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__469__A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high_inst/HI[324] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[70\]_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[6\]_B la_buf_enable\[6\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[3\] la_oenb_mprj[3] la_buf_enable\[3\]/B vssd vssd vccd vccd la_buf\[3\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__379__A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[34\] la_iena_mprj[34] mprj_logic_high_inst/HI[364] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[34\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[61\]_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[12\] la_oenb_mprj[12] la_buf_enable\[12\]/B vssd vssd vccd vccd la_buf\[12\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_10_1722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xpowergood_check vccd vdda2 mprj2_vdd_pwrgood/A mprj_vdd_pwrgood/A vdda1 vssd vssd
+ vssd vssd vdda1 mgmt_protect_hv
XFILLER_28_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[52\]_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] user_to_mprj_in_gates\[91\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[91\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[0\]_A _394_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[43\]_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[108\] _369_/Y mprj_logic_high_inst/HI[310] vssd vssd vccd
+ vccd la_oenb_core[108] sky130_fd_sc_hd__einvp_8
XFILLER_29_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[38\] _628_/Y mprj_logic_high_inst/HI[240] vssd vssd vccd
+ vccd la_oenb_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_38_2345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[34\]_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__572__A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[1\]_A _431_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y vssd vssd vccd vccd la_data_in_mprj[61]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[25\]_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__482__A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__657__A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[16\]_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__392__A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__567__A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_653_ la_oenb_mprj[63] vssd vssd vccd vccd _653_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[65\] _527_/Y la_buf\[65\]/TE vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__einvp_8
X_584_ la_data_out_mprj[122] vssd vssd vccd vccd _584_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[121\] _583_/Y la_buf\[121\]/TE vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[29\] _427_/Y mprj_adr_buf\[29\]/TE vssd vssd vccd vccd mprj_adr_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_32_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] user_to_mprj_in_gates\[54\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[54\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__477__A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__387__A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[54\]_A user_to_mprj_in_gates\[54\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[101\]_A_N la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_636_ la_oenb_mprj[46] vssd vssd vccd vccd _636_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[116\]_A_N la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_567_ la_data_out_mprj[105] vssd vssd vccd vccd _567_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_498_ la_data_out_mprj[36] vssd vssd vccd vccd _498_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y vssd vssd vccd vccd la_data_in_mprj[24]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[85\]_A _547_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[64\] la_iena_mprj[64] mprj_logic_high_inst/HI[394] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[64\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[2\] _592_/Y mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd la_oenb_core[2] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[20\] _610_/Y mprj_logic_high_inst/HI[222] vssd vssd vccd
+ vccd la_oenb_core[20] sky130_fd_sc_hd__einvp_8
X_421_ mprj_adr_o_core[23] vssd vssd vccd vccd _421_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[42\] la_oenb_mprj[42] la_buf_enable\[42\]/B vssd vssd vccd vccd la_buf\[42\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_352_ la_oenb_mprj[91] vssd vssd vccd vccd _352_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[94\]_B la_buf_enable\[94\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__580__A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[28\] _490_/Y la_buf\[28\]/TE vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__einvp_8
XFILLER_5_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_619_ la_oenb_mprj[29] vssd vssd vccd vccd _619_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[67\]_A _529_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] user_to_mprj_in_gates\[17\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[17\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[85\]_B la_buf_enable\[85\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__490__A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[76\]_B la_buf_enable\[76\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[68\] _329_/Y mprj_logic_high_inst/HI[270] vssd vssd vccd
+ vccd la_oenb_core[68] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[16\] _446_/Y mprj_dat_buf\[16\]/TE vssd vssd vccd vccd mprj_dat_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__575__A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_404_ mprj_adr_o_core[6] vssd vssd vccd vccd _404_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_335_ la_oenb_mprj[74] vssd vssd vccd vccd _335_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_B la_buf_enable\[67\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[11\] _409_/Y mprj_adr_buf\[11\]/TE vssd vssd vccd vccd mprj_adr_o_user[11]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[125] sky130_fd_sc_hd__inv_8
XFILLER_29_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y vssd vssd vccd vccd la_data_in_mprj[91]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__485__A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__395__A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[61\]_B mprj_logic_high_inst/HI[391] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[27\] la_iena_mprj[27] mprj_logic_high_inst/HI[357] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[27\]/B sky130_fd_sc_hd__and2_1
XFILLER_23_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[49\]_B la_buf_enable\[49\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_2159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[74\]_A_N la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[95\] _557_/Y la_buf\[95\]/TE vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[0\] la_iena_mprj[0] mprj_logic_high_inst/HI[330] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[0\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[110\] la_oenb_mprj[110] la_buf_enable\[110\]/B vssd vssd vccd vccd
+ la_buf\[110\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[89\]_A_N la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[52\]_B mprj_logic_high_inst/HI[382] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[12\]_A_N la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[9\]_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[27\]_A_N la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] user_to_mprj_in_gates\[84\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[84\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[43\]_B mprj_logic_high_inst/HI[373] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[34\]_B mprj_logic_high_inst/HI[364] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_32_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[6\] _468_/Y la_buf\[6\]/TE vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__einvp_8
XFILLER_10_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[10\] _472_/Y la_buf\[10\]/TE vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_3_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[3\] _401_/Y mprj_adr_buf\[3\]/TE vssd vssd vccd vccd mprj_adr_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[20\]_A _418_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y vssd vssd vccd vccd la_data_in_mprj[54]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[25\]_B mprj_logic_high_inst/HI[355] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high_inst/HI[213] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] user_to_mprj_in_gates\[110\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[110\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_27_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[16\]_B mprj_logic_high_inst/HI[346] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[94\] la_iena_mprj[94] mprj_logic_high_inst/HI[424] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[94\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[120\] _381_/Y mprj_logic_high_inst/HI[322] vssd vssd vccd
+ vccd la_oenb_core[120] sky130_fd_sc_hd__einvp_8
XFILLER_1_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[1\] _395_/Y mprj_sel_buf\[1\]/TE vssd vssd vccd vccd mprj_sel_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_27_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[50\] _640_/Y mprj_logic_high_inst/HI[252] vssd vssd vccd
+ vccd la_oenb_core[50] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[72\] la_oenb_mprj[72] la_buf_enable\[72\]/B vssd vssd vccd vccd la_buf\[72\]/TE
+ sky130_fd_sc_hd__and2b_1
X_652_ la_oenb_mprj[62] vssd vssd vccd vccd _652_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_583_ la_data_out_mprj[121] vssd vssd vccd vccd _583_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__583__A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[58\] _520_/Y la_buf\[58\]/TE vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__einvp_8
XFILLER_38_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[34\]_TE mprj_logic_high_inst/HI[236] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[114\] _576_/Y la_buf\[114\]/TE vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_10_1350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] user_to_mprj_in_gates\[47\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[47\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__493__A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] user_to_mprj_in_gates\[9\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[9\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_2334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[72\]_TE la_buf\[72\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[98\] _359_/Y mprj_logic_high_inst/HI[300] vssd vssd vccd
+ vccd la_oenb_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_29_1419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__578__A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_635_ la_oenb_mprj[45] vssd vssd vccd vccd _635_/Y sky130_fd_sc_hd__inv_2
X_566_ la_data_out_mprj[104] vssd vssd vccd vccd _566_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_497_ la_data_out_mprj[35] vssd vssd vccd vccd _497_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[0\]_TE mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y vssd vssd vccd vccd la_data_in_mprj[17]
+ sky130_fd_sc_hd__inv_8
XFILLER_5_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__488__A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[15\]_A _445_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__398__A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[57\] la_iena_mprj[57] mprj_logic_high_inst/HI[387] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[57\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_420_ mprj_adr_o_core[22] vssd vssd vccd vccd _420_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[13\] _603_/Y mprj_logic_high_inst/HI[215] vssd vssd vccd
+ vccd la_oenb_core[13] sky130_fd_sc_hd__einvp_8
X_351_ la_oenb_mprj[90] vssd vssd vccd vccd _351_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[35\] la_oenb_mprj[35] la_buf_enable\[35\]/B vssd vssd vccd vccd la_buf\[35\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y vssd vssd vccd vccd la_data_in_mprj[9]
+ sky130_fd_sc_hd__inv_8
XFILLER_35_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_618_ la_oenb_mprj[28] vssd vssd vccd vccd _618_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_549_ la_data_out_mprj[87] vssd vssd vccd vccd _549_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_A_N la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[115\]_A_N la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_403_ mprj_adr_o_core[5] vssd vssd vccd vccd _403_/Y sky130_fd_sc_hd__inv_2
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[40\] _502_/Y la_buf\[40\]/TE vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__einvp_8
X_334_ la_oenb_mprj[73] vssd vssd vccd vccd _334_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__591__A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[112\] la_iena_mprj[112] mprj_logic_high_inst/HI[442] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[112\]/B sky130_fd_sc_hd__and2_1
XFILLER_15_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[118] sky130_fd_sc_hd__inv_8
XFILLER_2_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y vssd vssd vccd vccd la_data_in_mprj[84]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_2317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[9\]_A _407_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[80\] _341_/Y mprj_logic_high_inst/HI[282] vssd vssd vccd
+ vccd la_oenb_core[80] sky130_fd_sc_hd__einvp_8
XFILLER_3_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__586__A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[88\] _550_/Y la_buf\[88\]/TE vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[103\] la_oenb_mprj[103] la_buf_enable\[103\]/B vssd vssd vccd vccd
+ la_buf\[103\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_19_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[9\]_B mprj_logic_high_inst/HI[339] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] user_to_mprj_in_gates\[77\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[77\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__496__A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high_inst/HI[292] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y vssd vssd vccd vccd la_data_in_mprj[47]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] user_to_mprj_in_gates\[103\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[103\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[73\]_A_N la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[88\]_A_N la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[87\] la_iena_mprj[87] mprj_logic_high_inst/HI[417] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[87\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[113\] _374_/Y mprj_logic_high_inst/HI[315] vssd vssd vccd
+ vccd la_oenb_core[113] sky130_fd_sc_hd__einvp_8
Xmprj_clk2_buf _390_/Y mprj_clk2_buf/TE vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__einvp_8
XFILLER_27_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[11\]_A_N la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[43\] _633_/Y mprj_logic_high_inst/HI[245] vssd vssd vccd
+ vccd la_oenb_core[43] sky130_fd_sc_hd__einvp_8
X_651_ la_oenb_mprj[61] vssd vssd vccd vccd _651_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[65\] la_oenb_mprj[65] la_buf_enable\[65\]/B vssd vssd vccd vccd la_buf\[65\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_irq_buffers\[1\] user_irq_gates\[1\]/Y vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__inv_8
X_582_ la_data_out_mprj[120] vssd vssd vccd vccd _582_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[26\]_A_N la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2188 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[107\] _569_/Y la_buf\[107\]/TE vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[100] sky130_fd_sc_hd__inv_8
XFILLER_0_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[120\]_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high_inst/HI[304] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[111\]_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1095 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_634_ la_oenb_mprj[44] vssd vssd vccd vccd _634_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__594__A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[70\] _532_/Y la_buf\[70\]/TE vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__einvp_8
XFILLER_17_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_565_ la_data_out_mprj[103] vssd vssd vccd vccd _565_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[102\]_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_496_ la_data_out_mprj[34] vssd vssd vccd vccd _496_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high_inst/HI[327] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[91\]_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_350_ la_oenb_mprj[89] vssd vssd vccd vccd _350_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[28\] la_oenb_mprj[28] la_buf_enable\[28\]/B vssd vssd vccd vccd la_buf\[28\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_6_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__589__A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[82\]_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_617_ la_oenb_mprj[27] vssd vssd vccd vccd _617_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_548_ la_data_out_mprj[86] vssd vssd vccd vccd _548_/Y sky130_fd_sc_hd__inv_2
X_479_ la_data_out_mprj[17] vssd vssd vccd vccd _479_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high_inst/HI[249] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__499__A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[73\]_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[9\]_B la_buf_enable\[9\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[64\]_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_402_ mprj_adr_o_core[4] vssd vssd vccd vccd _402_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_333_ la_oenb_mprj[72] vssd vssd vccd vccd _333_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[33\] _495_/Y la_buf\[33\]/TE vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[105\] la_iena_mprj[105] mprj_logic_high_inst/HI[435] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[105\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y vssd vssd vccd vccd la_data_in_mprj[77]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[55\]_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] user_to_mprj_in_gates\[22\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[22\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_sel_buf\[3\]_A _397_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[46\]_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[73\] _334_/Y mprj_logic_high_inst/HI[275] vssd vssd vccd
+ vccd la_oenb_core[73] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[95\] la_oenb_mprj[95] la_buf_enable\[95\]/B vssd vssd vccd vccd la_buf\[95\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[21\] _451_/Y mprj_dat_buf\[21\]/TE vssd vssd vccd vccd mprj_dat_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[37\]_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1848 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[28\]_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[114\]_A_N la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[1\] la_oenb_mprj[1] la_buf_enable\[1\]/B vssd vssd vccd vccd la_buf\[1\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_2150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[19\]_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[32\] la_iena_mprj[32] mprj_logic_high_inst/HI[362] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[32\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[10\] la_oenb_mprj[10] la_buf_enable\[10\]/B vssd vssd vccd vccd la_buf\[10\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__597__A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[111\]_A _573_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _367_/Y mprj_logic_high_inst/HI[308] vssd vssd vccd
+ vccd la_oenb_core[106] sky130_fd_sc_hd__einvp_8
XFILLER_5_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_650_ la_oenb_mprj[60] vssd vssd vccd vccd _650_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[36\] _626_/Y mprj_logic_high_inst/HI[238] vssd vssd vccd
+ vccd la_oenb_core[36] sky130_fd_sc_hd__einvp_8
X_581_ la_data_out_mprj[119] vssd vssd vccd vccd _581_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[58\] la_oenb_mprj[58] la_buf_enable\[58\]/B vssd vssd vccd vccd la_buf\[58\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_17_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high_inst/HI[282] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[120\]_B mprj_logic_high_inst/HI[450] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[21\]_A _483_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[88\]_A _550_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[111\]_B mprj_logic_high_inst/HI[441] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[12\]_A _474_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[30\]_B la_buf_enable\[30\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_633_ la_oenb_mprj[43] vssd vssd vccd vccd _633_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[79\]_A _541_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[63\] _525_/Y la_buf\[63\]/TE vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__einvp_8
X_564_ la_data_out_mprj[102] vssd vssd vccd vccd _564_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[102\]_B mprj_logic_high_inst/HI[432] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_495_ la_data_out_mprj[33] vssd vssd vccd vccd _495_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[97\]_B la_buf_enable\[97\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[27\] _425_/Y mprj_adr_buf\[27\]/TE vssd vssd vccd vccd mprj_adr_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_23_2200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[21\]_B la_buf_enable\[21\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[72\]_A_N la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] user_to_mprj_in_gates\[52\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[52\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[87\]_A_N la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[88\]_B la_buf_enable\[88\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[10\]_A_N la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[25\]_A_N la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[12\]_B la_buf_enable\[12\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[91\]_B mprj_logic_high_inst/HI[421] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[79\]_B la_buf_enable\[79\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[81\]_A _342_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[126\] la_oenb_mprj[126] la_buf_enable\[126\]/B vssd vssd vccd vccd
+ la_buf\[126\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_24_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_616_ la_oenb_mprj[26] vssd vssd vccd vccd _616_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_547_ la_data_out_mprj[85] vssd vssd vccd vccd _547_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_478_ la_data_out_mprj[16] vssd vssd vccd vccd _478_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y vssd vssd vccd vccd la_data_in_mprj[22]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[62\] la_iena_mprj[62] mprj_logic_high_inst/HI[392] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[62\]/B sky130_fd_sc_hd__and2_1
XFILLER_18_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[64\]_B mprj_logic_high_inst/HI[394] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[0\] _590_/Y mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd la_oenb_core[0] sky130_fd_sc_hd__einvp_8
X_401_ mprj_adr_o_core[3] vssd vssd vccd vccd _401_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[40\] la_oenb_mprj[40] la_buf_enable\[40\]/B vssd vssd vccd vccd la_buf\[40\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_332_ la_oenb_mprj[71] vssd vssd vccd vccd _332_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high_inst/HI[317] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[26\] _488_/Y la_buf\[26\]/TE vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_6_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[55\]_B mprj_logic_high_inst/HI[385] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] user_to_mprj_in_gates\[15\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[15\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high_inst/HI[216] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] user_to_mprj_in_gates\[126\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[126\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[46\]_B mprj_logic_high_inst/HI[376] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[66\] _656_/Y mprj_logic_high_inst/HI[268] vssd vssd vccd
+ vccd la_oenb_core[66] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[88\] la_oenb_mprj[88] la_buf_enable\[88\]/B vssd vssd vccd vccd la_buf\[88\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[14\] _444_/Y mprj_dat_buf\[14\]/TE vssd vssd vccd vccd mprj_dat_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[37\]_B mprj_logic_high_inst/HI[367] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[37\]_TE mprj_logic_high_inst/HI[239] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_843 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[123] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_adr_buf\[23\]_A _421_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[28\]_B mprj_logic_high_inst/HI[358] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[75\]_TE la_buf\[75\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[14\]_A _412_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[19\]_B mprj_logic_high_inst/HI[349] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[25\] la_iena_mprj[25] mprj_logic_high_inst/HI[355] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[25\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[93\] _555_/Y la_buf\[93\]/TE vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_1_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] user_to_mprj_in_gates\[82\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[82\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_580_ la_data_out_mprj[118] vssd vssd vccd vccd _580_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[29\] _619_/Y mprj_logic_high_inst/HI[231] vssd vssd vccd
+ vccd la_oenb_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_31_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[4\] _466_/Y la_buf\[4\]/TE vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__einvp_8
XFILLER_10_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[113\]_A_N la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__401__A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[1\] _399_/Y mprj_adr_buf\[1\]/TE vssd vssd vccd vccd mprj_adr_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_23_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y vssd vssd vccd vccd la_data_in_mprj[52]
+ sky130_fd_sc_hd__inv_8
XFILLER_23_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_A _448_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[100\]_TE la_buf\[100\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[92\] la_iena_mprj[92] mprj_logic_high_inst/HI[422] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[92\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[70\] la_oenb_mprj[70] la_buf_enable\[70\]/B vssd vssd vccd vccd la_buf\[70\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_632_ la_oenb_mprj[42] vssd vssd vccd vccd _632_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_563_ la_data_out_mprj[101] vssd vssd vccd vccd _563_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[56\] _518_/Y la_buf\[56\]/TE vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__einvp_8
X_494_ la_data_out_mprj[32] vssd vssd vccd vccd _494_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[112\] _574_/Y la_buf\[112\]/TE vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__einvp_8
XFILLER_29_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[120\]_B la_buf_enable\[120\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] user_to_mprj_in_gates\[45\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[45\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[123\]_TE la_buf\[123\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] user_to_mprj_in_gates\[7\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[7\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[111\]_B la_buf_enable\[111\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[96\] _357_/Y mprj_logic_high_inst/HI[298] vssd vssd vccd
+ vccd la_oenb_core[96] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[9\] la_iena_mprj[9] mprj_logic_high_inst/HI[339] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[9\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_1820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[119\] la_oenb_mprj[119] la_buf_enable\[119\]/B vssd vssd vccd vccd
+ la_buf\[119\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_615_ la_oenb_mprj[25] vssd vssd vccd vccd _615_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[102\]_B la_buf_enable\[102\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_546_ la_data_out_mprj[84] vssd vssd vccd vccd _546_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_477_ la_data_out_mprj[15] vssd vssd vccd vccd _477_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y vssd vssd vccd vccd la_data_in_mprj[15]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high_inst/HI[295] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_pwrgood mprj2_pwrgood/A vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_8_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[55\] la_iena_mprj[55] mprj_logic_high_inst/HI[385] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[55\]/B sky130_fd_sc_hd__and2_1
XFILLER_18_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_400_ mprj_adr_o_core[2] vssd vssd vccd vccd _400_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[11\] _601_/Y mprj_logic_high_inst/HI[213] vssd vssd vccd
+ vccd la_oenb_core[11] sky130_fd_sc_hd__einvp_8
X_331_ la_oenb_mprj[70] vssd vssd vccd vccd _331_/Y sky130_fd_sc_hd__inv_2
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y vssd vssd vccd vccd la_data_in_mprj[7]
+ sky130_fd_sc_hd__inv_8
Xla_buf_enable\[33\] la_oenb_mprj[33] la_buf_enable\[33\]/B vssd vssd vccd vccd la_buf\[33\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[71\]_A_N la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[19\] _481_/Y la_buf\[19\]/TE vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_6_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[86\]_A_N la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[24\]_A_N la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_529_ la_data_out_mprj[67] vssd vssd vccd vccd _529_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[39\]_A_N la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_vdd_pwrgood_A mprj_vdd_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] user_to_mprj_in_gates\[119\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[119\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[59\] _649_/Y mprj_logic_high_inst/HI[261] vssd vssd vccd
+ vccd la_oenb_core[59] sky130_fd_sc_hd__einvp_8
XFILLER_1_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[110\] la_iena_mprj[110] mprj_logic_high_inst/HI[440] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[110\]/B sky130_fd_sc_hd__and2_1
XFILLER_15_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__404__A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[116] sky130_fd_sc_hd__inv_8
XFILLER_2_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y vssd vssd vccd vccd la_data_in_mprj[82]
+ sky130_fd_sc_hd__inv_8
XFILLER_38_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[105\]_TE mprj_logic_high_inst/HI[307] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[18\] la_iena_mprj[18] mprj_logic_high_inst/HI[348] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[18\]/B sky130_fd_sc_hd__and2_1
XFILLER_12_637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[86\] _548_/Y la_buf\[86\]/TE vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[101\] la_oenb_mprj[101] la_buf_enable\[101\]/B vssd vssd vccd vccd
+ la_buf\[101\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_5_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] user_to_mprj_in_gates\[75\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[75\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[123\]_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2203 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high_inst/HI[229] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[114\]_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_2147 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_427 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_ena_buf\[1\] user_irq_ena[1] user_irq_ena_buf\[1\]/B vssd vssd vccd vccd
+ user_irq_gates\[1\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[105\]_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y vssd vssd vccd vccd la_data_in_mprj[45]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_950 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] user_to_mprj_in_gates\[101\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[101\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_21_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__502__A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[85\] la_iena_mprj[85] mprj_logic_high_inst/HI[415] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[85\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[111\] _372_/Y mprj_logic_high_inst/HI[313] vssd vssd vccd
+ vccd la_oenb_core[111] sky130_fd_sc_hd__einvp_8
XFILLER_0_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[94\]_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[41\] _631_/Y mprj_logic_high_inst/HI[243] vssd vssd vccd
+ vccd la_oenb_core[41] sky130_fd_sc_hd__einvp_8
X_631_ la_oenb_mprj[41] vssd vssd vccd vccd _631_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[63\] la_oenb_mprj[63] la_buf_enable\[63\]/B vssd vssd vccd vccd la_buf\[63\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_562_ la_data_out_mprj[100] vssd vssd vccd vccd _562_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_493_ la_data_out_mprj[31] vssd vssd vccd vccd _493_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[49\] _511_/Y la_buf\[49\]/TE vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_9_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__412__A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[105\] _567_/Y la_buf\[105\]/TE vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[85\]_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] user_to_mprj_in_gates\[38\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[38\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[76\]_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[112\]_A_N la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[127\]_A_N la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[89\] _350_/Y mprj_logic_high_inst/HI[291] vssd vssd vccd
+ vccd la_oenb_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_1_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[67\]_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_614_ la_oenb_mprj[24] vssd vssd vccd vccd _614_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_545_ la_data_out_mprj[83] vssd vssd vccd vccd _545_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__407__A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_476_ la_data_out_mprj[14] vssd vssd vccd vccd _476_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[58\]_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2087 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[49\]_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[48\] la_iena_mprj[48] mprj_logic_high_inst/HI[378] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[48\]/B sky130_fd_sc_hd__and2_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_330_ la_oenb_mprj[69] vssd vssd vccd vccd _330_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[26\] la_oenb_mprj[26] la_buf_enable\[26\]/B vssd vssd vccd vccd la_buf\[26\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_17_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[28\]_TE mprj_adr_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[7\]_A _437_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_528_ la_data_out_mprj[66] vssd vssd vccd vccd _528_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_370 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_459_ mprj_dat_o_core[29] vssd vssd vccd vccd _459_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__600__A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__510__A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_646 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[31\] _493_/Y la_buf\[31\]/TE vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[103\] la_iena_mprj[103] mprj_logic_high_inst/HI[433] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[103\]/B sky130_fd_sc_hd__and2_1
XFILLER_7_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[110\]_B user_to_mprj_in_gates\[110\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high_inst/HI[285] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__420__A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[109] sky130_fd_sc_hd__inv_8
XFILLER_20_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y vssd vssd vccd vccd la_data_in_mprj[75]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] user_to_mprj_in_gates\[20\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[20\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_34_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[125\]_A user_to_mprj_in_gates\[125\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__330__A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[8\] _438_/Y mprj_dat_buf\[8\]/TE vssd vssd vccd vccd mprj_dat_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[70\]_A_N la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[85\]_A_N la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__505__A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[69\]_A user_to_mprj_in_gates\[69\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[23\]_A_N la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[71\] _332_/Y mprj_logic_high_inst/HI[273] vssd vssd vccd
+ vccd la_oenb_core[71] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[93\] la_oenb_mprj[93] la_buf_enable\[93\]/B vssd vssd vccd vccd la_buf\[93\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_23_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[38\]_A_N la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[79\] _541_/Y la_buf\[79\]/TE vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_31_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__415__A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] user_to_mprj_in_gates\[68\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[68\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[123\]_B mprj_logic_high_inst/HI[453] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_18_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[24\]_A _486_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[42\]_B la_buf_enable\[42\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[114\]_B mprj_logic_high_inst/HI[444] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[30\] la_iena_mprj[30] mprj_logic_high_inst/HI[360] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[30\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_2159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1311 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[15\]_A _477_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[33\]_B la_buf_enable\[33\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[2\]_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[105\]_B mprj_logic_high_inst/HI[435] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y vssd vssd vccd vccd la_data_in_mprj[38]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf_enable\[24\]_B la_buf_enable\[24\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[15\]_B la_buf_enable\[15\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[78\] la_iena_mprj[78] mprj_logic_high_inst/HI[408] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[78\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[94\]_B mprj_logic_high_inst/HI[424] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[104\] _365_/Y mprj_logic_high_inst/HI[306] vssd vssd vccd
+ vccd la_oenb_core[104] sky130_fd_sc_hd__einvp_8
X_630_ la_oenb_mprj[40] vssd vssd vccd vccd _630_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[34\] _624_/Y mprj_logic_high_inst/HI[236] vssd vssd vccd
+ vccd la_oenb_core[34] sky130_fd_sc_hd__einvp_8
X_561_ la_data_out_mprj[99] vssd vssd vccd vccd _561_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[56\] la_oenb_mprj[56] la_buf_enable\[56\]/B vssd vssd vccd vccd la_buf\[56\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_492_ la_data_out_mprj[30] vssd vssd vccd vccd _492_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_715 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high_inst/HI[320] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[85\]_B mprj_logic_high_inst/HI[415] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[17\]_TE mprj_logic_high_inst/HI[219] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__603__A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_2219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__513__A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[67\]_B mprj_logic_high_inst/HI[397] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_29_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_613_ la_oenb_mprj[23] vssd vssd vccd vccd _613_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_1938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[61\] _523_/Y la_buf\[61\]/TE vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__einvp_8
X_544_ la_data_out_mprj[82] vssd vssd vccd vccd _544_/Y sky130_fd_sc_hd__inv_2
X_475_ la_data_out_mprj[13] vssd vssd vccd vccd _475_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__423__A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[25\] _423_/Y mprj_adr_buf\[25\]/TE vssd vssd vccd vccd mprj_adr_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[58\]_B mprj_logic_high_inst/HI[388] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2099 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1415 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] user_to_mprj_in_gates\[50\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[50\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__333__A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[49\]_B mprj_logic_high_inst/HI[379] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__508__A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[19\] la_oenb_mprj[19] la_buf_enable\[19\]/B vssd vssd vccd vccd la_buf\[19\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_irq_gates\[2\] user_irq_core[2] user_irq_gates\[2\]/B vssd vssd vccd vccd user_irq_gates\[2\]/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[124\] la_oenb_mprj[124] la_buf_enable\[124\]/B vssd vssd vccd vccd
+ la_buf\[124\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_18_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[27\]_TE mprj_dat_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__418__A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_527_ la_data_out_mprj[65] vssd vssd vccd vccd _527_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[6\]_TE mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_458_ mprj_dat_o_core[28] vssd vssd vccd vccd _458_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_389_ caravel_clk vssd vssd vccd vccd _389_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y vssd vssd vccd vccd la_data_in_mprj[20]
+ sky130_fd_sc_hd__inv_8
XFILLER_31_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] user_to_mprj_in_gates\[98\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[98\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[26\]_A _424_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[111\]_A_N la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[126\]_A_N la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[3\]_A _593_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[60\] la_iena_mprj[60] mprj_logic_high_inst/HI[390] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[60\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[24\] _486_/Y la_buf\[24\]/TE vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__einvp_8
XFILLER_6_323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y vssd vssd vccd vccd la_data_in_mprj[68]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] user_to_mprj_in_gates\[13\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[13\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__611__A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] user_to_mprj_in_gates\[124\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[124\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__521__A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[64\] _654_/Y mprj_logic_high_inst/HI[266] vssd vssd vccd
+ vccd la_oenb_core[64] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[86\] la_oenb_mprj[86] la_buf_enable\[86\]/B vssd vssd vccd vccd la_buf\[86\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[12\] _442_/Y mprj_dat_buf\[12\]/TE vssd vssd vccd vccd mprj_dat_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XFILLER_28_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[50\]_TE mprj_logic_high_inst/HI[252] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__431__A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[121] sky130_fd_sc_hd__inv_8
XFILLER_26_2234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__606__A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[2\]_A _400_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__341__A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[73\]_TE mprj_logic_high_inst/HI[275] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[23\] la_iena_mprj[23] mprj_logic_high_inst/HI[353] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[23\]/B sky130_fd_sc_hd__and2_1
XANTENNA__516__A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[2\]_B mprj_logic_high_inst/HI[332] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[91\] _553_/Y la_buf\[91\]/TE vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_5_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__426__A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] user_to_mprj_in_gates\[80\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[80\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[84\]_A_N la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high_inst/HI[298] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[123\]_B la_buf_enable\[123\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[99\]_A_N la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_A_N la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__336__A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[37\]_A_N la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[114\]_B la_buf_enable\[114\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_560_ la_data_out_mprj[98] vssd vssd vccd vccd _560_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[27\] _617_/Y mprj_logic_high_inst/HI[229] vssd vssd vccd
+ vccd la_oenb_core[27] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[9\] _599_/Y mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd la_oenb_core[9] sky130_fd_sc_hd__einvp_8
X_491_ la_data_out_mprj[29] vssd vssd vccd vccd _491_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[49\] la_oenb_mprj[49] la_buf_enable\[49\]/B vssd vssd vccd vccd la_buf\[49\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[2\] _464_/Y la_buf\[2\]/TE vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__einvp_8
XFILLER_5_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_660 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[8\]_A _470_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[105\]_B la_buf_enable\[105\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y vssd vssd vccd vccd la_data_in_mprj[50]
+ sky130_fd_sc_hd__inv_8
XFILLER_35_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_737 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[90\] la_iena_mprj[90] mprj_logic_high_inst/HI[420] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[90\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_612_ la_oenb_mprj[22] vssd vssd vccd vccd _612_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_543_ la_data_out_mprj[81] vssd vssd vccd vccd _543_/Y sky130_fd_sc_hd__inv_2
X_474_ la_data_out_mprj[12] vssd vssd vccd vccd _474_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[54\] _516_/Y la_buf\[54\]/TE vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[126\] la_iena_mprj[126] mprj_logic_high_inst/HI[456] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[126\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[110\] _572_/Y la_buf\[110\]/TE vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[18\] _416_/Y mprj_adr_buf\[18\]/TE vssd vssd vccd vccd mprj_adr_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y vssd vssd vccd vccd la_data_in_mprj[98]
+ sky130_fd_sc_hd__inv_8
XFILLER_23_2023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] user_to_mprj_in_gates\[43\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[43\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_35_199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__614__A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] user_to_mprj_in_gates\[5\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[5\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_2039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[108\]_TE mprj_logic_high_inst/HI[310] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__524__A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[94\] _355_/Y mprj_logic_high_inst/HI[296] vssd vssd vccd
+ vccd la_oenb_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_1_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[7\] la_iena_mprj[7] mprj_logic_high_inst/HI[337] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[7\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[117\] la_oenb_mprj[117] la_buf_enable\[117\]/B vssd vssd vccd vccd
+ la_buf\[117\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_24_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_526_ la_data_out_mprj[64] vssd vssd vccd vccd _526_/Y sky130_fd_sc_hd__inv_2
X_457_ mprj_dat_o_core[27] vssd vssd vccd vccd _457_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_388_ la_oenb_mprj[127] vssd vssd vccd vccd _388_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__434__A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y vssd vssd vccd vccd la_data_in_mprj[13]
+ sky130_fd_sc_hd__inv_8
XFILLER_5_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__609__A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__344__A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[53\] la_iena_mprj[53] mprj_logic_high_inst/HI[383] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[53\]/B sky130_fd_sc_hd__and2_1
XANTENNA__519__A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y vssd vssd vccd vccd la_data_in_mprj[5]
+ sky130_fd_sc_hd__inv_8
Xla_buf_enable\[31\] la_oenb_mprj[31] la_buf_enable\[31\]/B vssd vssd vccd vccd la_buf\[31\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_19_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[17\] _479_/Y la_buf\[17\]/TE vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__einvp_8
XFILLER_6_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__429__A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_509_ la_data_out_mprj[47] vssd vssd vccd vccd _509_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_128 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[2\]_B la_buf_enable\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[126\]_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] user_to_mprj_in_gates\[117\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[117\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__339__A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[127\] _388_/Y mprj_logic_high_inst/HI[329] vssd vssd vccd
+ vccd la_oenb_core[127] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[57\] _647_/Y mprj_logic_high_inst/HI[259] vssd vssd vccd
+ vccd la_oenb_core[57] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[79\] la_oenb_mprj[79] la_buf_enable\[79\]/B vssd vssd vccd vccd la_buf\[79\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[117\]_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_A_N la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[125\]_A_N la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[114] sky130_fd_sc_hd__inv_8
XFILLER_6_2318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y vssd vssd vccd vccd la_data_in_mprj[80]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[108\]_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__622__A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1976 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[16\] la_iena_mprj[16] mprj_logic_high_inst/HI[346] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[16\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[30\]_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__532__A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[97\]_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[84\] _546_/Y la_buf\[84\]/TE vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_1_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__442__A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[88\]_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] user_to_mprj_in_gates\[73\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[73\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__617__A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[12\]_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__352__A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[79\]_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high_inst/HI[242] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__527__A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_490_ la_data_out_mprj[28] vssd vssd vccd vccd _490_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1745 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__437__A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y vssd vssd vccd vccd la_data_in_mprj[43]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__347__A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_749 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[83\] la_iena_mprj[83] mprj_logic_high_inst/HI[413] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[83\]/B sky130_fd_sc_hd__and2_1
XFILLER_7_1019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[50\]_A user_to_mprj_in_gates\[50\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_611_ la_oenb_mprj[21] vssd vssd vccd vccd _611_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[61\] la_oenb_mprj[61] la_buf_enable\[61\]/B vssd vssd vccd vccd la_buf\[61\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_542_ la_data_out_mprj[80] vssd vssd vccd vccd _542_/Y sky130_fd_sc_hd__inv_2
X_473_ la_data_out_mprj[11] vssd vssd vccd vccd _473_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[47\] _509_/Y la_buf\[47\]/TE vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__einvp_8
XFILLER_13_565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[83\]_A_N la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[119\] la_iena_mprj[119] mprj_logic_high_inst/HI[449] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[119\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[90\]_A _552_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high_inst/HI[288] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[98\]_A_N la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[103\] _565_/Y la_buf\[103\]/TE vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__einvp_8
XFILLER_29_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[21\]_A_N la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_2035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[36\]_A_N la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] user_to_mprj_in_gates\[36\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[36\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[81\]_A _543_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__630__A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[72\]_A _534_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[90\]_B la_buf_enable\[90\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__540__A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[87\] _348_/Y mprj_logic_high_inst/HI[289] vssd vssd vccd
+ vccd la_oenb_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_1_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_525_ la_data_out_mprj[63] vssd vssd vccd vccd _525_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[126\]_A _588_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_456_ mprj_dat_o_core[26] vssd vssd vccd vccd _456_/Y sky130_fd_sc_hd__inv_2
X_387_ la_oenb_mprj[126] vssd vssd vccd vccd _387_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[113\]_B user_to_mprj_in_gates\[113\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[63\]_A _525_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[30\] _428_/Y mprj_adr_buf\[30\]/TE vssd vssd vccd vccd mprj_adr_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[81\]_B la_buf_enable\[81\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__450__A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[117\]_A _579_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__625__A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[54\]_A _516_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[72\]_B la_buf_enable\[72\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__360__A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_stb_buf_A _392_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[46\] la_iena_mprj[46] mprj_logic_high_inst/HI[376] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[46\]/B sky130_fd_sc_hd__and2_1
XFILLER_21_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__535__A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[24\] la_oenb_mprj[24] la_buf_enable\[24\]/B vssd vssd vccd vccd la_buf\[24\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_508_ la_data_out_mprj[46] vssd vssd vccd vccd _508_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__445__A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_439_ mprj_dat_o_core[9] vssd vssd vccd vccd _439_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[54\]_B la_buf_enable\[54\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[126\]_B mprj_logic_high_inst/HI[456] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__355__A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[27\]_A _489_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[45\]_B la_buf_enable\[45\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[117\]_B mprj_logic_high_inst/HI[447] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[18\]_A _480_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[101\] la_iena_mprj[101] mprj_logic_high_inst/HI[431] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[101\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[36\]_B la_buf_enable\[36\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[5\]_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[107] sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[108\]_B mprj_logic_high_inst/HI[438] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y vssd vssd vccd vccd la_data_in_mprj[73]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[27\]_B la_buf_enable\[27\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _436_/Y mprj_dat_buf\[6\]/TE vssd vssd vccd vccd mprj_dat_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[30\]_B mprj_logic_high_inst/HI[360] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[18\]_B la_buf_enable\[18\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[91\] la_oenb_mprj[91] la_buf_enable\[91\]/B vssd vssd vccd vccd la_buf\[91\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[97\]_B mprj_logic_high_inst/HI[427] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1916 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[58\]_TE la_buf\[58\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[77\] _539_/Y la_buf\[77\]/TE vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__einvp_8
XFILLER_38_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_B mprj_logic_high_inst/HI[351] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[88\]_B mprj_logic_high_inst/HI[418] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] user_to_mprj_in_gates\[66\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[66\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[12\]_B mprj_logic_high_inst/HI[342] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__633__A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[124\]_A_N la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__543__A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y vssd vssd vccd vccd la_data_in_mprj[36]
+ sky130_fd_sc_hd__inv_8
XANTENNA__453__A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__628__A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__363__A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[76\] la_iena_mprj[76] mprj_logic_high_inst/HI[406] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[76\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[102\] _363_/Y mprj_logic_high_inst/HI[304] vssd vssd vccd
+ vccd la_oenb_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_22_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_610_ la_oenb_mprj[20] vssd vssd vccd vccd _610_/Y sky130_fd_sc_hd__inv_2
XANTENNA__538__A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[32\] _622_/Y mprj_logic_high_inst/HI[234] vssd vssd vccd
+ vccd la_oenb_core[32] sky130_fd_sc_hd__einvp_8
X_541_ la_data_out_mprj[79] vssd vssd vccd vccd _541_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[54\] la_oenb_mprj[54] la_buf_enable\[54\]/B vssd vssd vccd vccd la_buf\[54\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_17_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_472_ la_data_out_mprj[10] vssd vssd vccd vccd _472_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[20\]_A _450_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_2047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__448__A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_820 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] user_to_mprj_in_gates\[29\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[29\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high_inst/HI[232] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[29\]_A _427_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__358__A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[6\]_A _596_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[28\] _458_/Y mprj_dat_buf\[28\]/TE vssd vssd vccd vccd mprj_dat_o_user[28]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_524_ la_data_out_mprj[62] vssd vssd vccd vccd _524_/Y sky130_fd_sc_hd__inv_2
X_455_ mprj_dat_o_core[25] vssd vssd vccd vccd _455_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_386_ la_oenb_mprj[125] vssd vssd vccd vccd _386_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[23\] _421_/Y mprj_adr_buf\[23\]/TE vssd vssd vccd vccd mprj_adr_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[9\]_TE mprj_dat_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[8\] la_oenb_mprj[8] la_buf_enable\[8\]/B vssd vssd vccd vccd la_buf\[8\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__641__A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[82\]_A_N la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[76\]_TE mprj_logic_high_inst/HI[278] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[39\] la_iena_mprj[39] mprj_logic_high_inst/HI[369] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[39\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[97\]_A_N la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[20\]_A_N la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[17\] la_oenb_mprj[17] la_buf_enable\[17\]/B vssd vssd vccd vccd la_buf\[17\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_6_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1957 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__551__A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[35\]_A_N la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_gates\[0\] user_irq_core[0] user_irq_gates\[0\]/B vssd vssd vccd vccd user_irq_gates\[0\]/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_2_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[122\] la_oenb_mprj[122] la_buf_enable\[122\]/B vssd vssd vccd vccd
+ la_buf\[122\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_24_2153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_507_ la_data_out_mprj[45] vssd vssd vccd vccd _507_/Y sky130_fd_sc_hd__inv_2
X_438_ mprj_dat_o_core[8] vssd vssd vccd vccd _438_/Y sky130_fd_sc_hd__inv_2
X_369_ la_oenb_mprj[108] vssd vssd vccd vccd _369_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__461__A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] user_to_mprj_in_gates\[96\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[96\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high_inst/HI[301] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__636__A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[5\]_A _403_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__371__A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__546__A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[22\] _484_/Y la_buf\[22\]/TE vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__einvp_8
XFILLER_6_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[5\]_B mprj_logic_high_inst/HI[335] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y vssd vssd vccd vccd la_data_in_mprj[66]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_stb_buf_TE mprj_stb_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__456__A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] user_to_mprj_in_gates\[11\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[11\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_1941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[126\]_B la_buf_enable\[126\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] user_to_mprj_in_gates\[122\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[122\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__366__A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[62\] _652_/Y mprj_logic_high_inst/HI[264] vssd vssd vccd
+ vccd la_oenb_core[62] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[84\] la_oenb_mprj[84] la_buf_enable\[84\]/B vssd vssd vccd vccd la_buf\[84\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[117\]_B la_buf_enable\[117\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[10\] _440_/Y mprj_dat_buf\[10\]/TE vssd vssd vccd vccd mprj_dat_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[126\] _588_/Y la_buf\[126\]/TE vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_6_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[108\]_B la_buf_enable\[108\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] user_to_mprj_in_gates\[59\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[59\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_19_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[21\] la_iena_mprj[21] mprj_logic_high_inst/HI[351] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[21\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y vssd vssd vccd vccd la_data_in_mprj[29]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__644__A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[48\]_TE la_buf\[48\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[69\] la_iena_mprj[69] mprj_logic_high_inst/HI[399] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[69\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_1600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_540_ la_data_out_mprj[78] vssd vssd vccd vccd _540_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[7\] _597_/Y mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd la_oenb_core[7] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[25\] _615_/Y mprj_logic_high_inst/HI[227] vssd vssd vccd
+ vccd la_oenb_core[25] sky130_fd_sc_hd__einvp_8
X_471_ la_data_out_mprj[9] vssd vssd vccd vccd _471_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[47\] la_oenb_mprj[47] la_buf_enable\[47\]/B vssd vssd vccd vccd la_buf\[47\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__554__A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[0\] _462_/Y la_buf\[0\]/TE vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__einvp_8
XFILLER_5_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__464__A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[123\]_A_N la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__639__A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__374__A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__549__A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_523_ la_data_out_mprj[61] vssd vssd vccd vccd _523_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_454_ mprj_dat_o_core[24] vssd vssd vccd vccd _454_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[52\] _514_/Y la_buf\[52\]/TE vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[124\] la_iena_mprj[124] mprj_logic_high_inst/HI[454] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[124\]/B sky130_fd_sc_hd__and2_1
X_385_ la_oenb_mprj[124] vssd vssd vccd vccd _385_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_2307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[16\] _414_/Y mprj_adr_buf\[16\]/TE vssd vssd vccd vccd mprj_adr_o_user[16]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y vssd vssd vccd vccd la_data_in_mprj[96]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__459__A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_rstn_buf caravel_rstn mprj_rstn_buf/TE vssd vssd vccd vccd user_reset sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] user_to_mprj_in_gates\[41\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[41\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[5\]_B la_buf_enable\[5\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] user_to_mprj_in_gates\[3\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[3\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__369__A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[121\]_TE mprj_logic_high_inst/HI[323] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[60\]_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[92\] _353_/Y mprj_logic_high_inst/HI[294] vssd vssd vccd
+ vccd la_oenb_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_2_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[5\] la_iena_mprj[5] mprj_logic_high_inst/HI[335] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[5\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_2165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[115\] la_oenb_mprj[115] la_buf_enable\[115\]/B vssd vssd vccd vccd
+ la_buf\[115\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[20\]_TE mprj_logic_high_inst/HI[222] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_506_ la_data_out_mprj[44] vssd vssd vccd vccd _506_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[51\]_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_437_ mprj_dat_o_core[7] vssd vssd vccd vccd _437_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_368_ la_oenb_mprj[107] vssd vssd vccd vccd _368_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y vssd vssd vccd vccd la_data_in_mprj[11]
+ sky130_fd_sc_hd__inv_8
XFILLER_5_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] user_to_mprj_in_gates\[89\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[89\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[42\]_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__652__A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[51\] la_iena_mprj[51] mprj_logic_high_inst/HI[381] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[51\]/B sky130_fd_sc_hd__and2_1
XFILLER_19_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_cyc_buf _391_/Y mprj_cyc_buf/TE vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__einvp_8
XFILLER_27_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[33\]_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_418 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y vssd vssd vccd vccd la_data_in_mprj[3]
+ sky130_fd_sc_hd__inv_8
XFILLER_30_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__562__A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[15\] _477_/Y la_buf\[15\]/TE vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[0\]_A _430_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_2205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[8\] _406_/Y mprj_adr_buf\[8\]/TE vssd vssd vccd vccd mprj_adr_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y vssd vssd vccd vccd la_data_in_mprj[59]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[24\]_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__472__A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[81\]_A_N la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[96\]_A_N la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] user_to_mprj_in_gates\[115\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[115\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__647__A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[34\]_A_N la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[15\]_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1786 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__382__A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[49\]_A_N la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[99\] la_iena_mprj[99] mprj_logic_high_inst/HI[429] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[99\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_1338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[30\]_TE mprj_dat_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[125\] _386_/Y mprj_logic_high_inst/HI[327] vssd vssd vccd
+ vccd la_oenb_core[125] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[55\] _645_/Y mprj_logic_high_inst/HI[257] vssd vssd vccd
+ vccd la_oenb_core[55] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[77\] la_oenb_mprj[77] la_buf_enable\[77\]/B vssd vssd vccd vccd la_buf\[77\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[2\]_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__557__A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high_inst/HI[291] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[119\] _581_/Y la_buf\[119\]/TE vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[112] sky130_fd_sc_hd__inv_8
XFILLER_6_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[71\]_A user_to_mprj_in_gates\[71\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__467__A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__377__A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[14\] la_iena_mprj[14] mprj_logic_high_inst/HI[344] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[14\]/B sky130_fd_sc_hd__and2_1
XFILLER_20_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[82\] _544_/Y la_buf\[82\]/TE vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__einvp_8
XFILLER_5_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] user_to_mprj_in_gates\[71\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[71\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_470_ la_data_out_mprj[8] vssd vssd vccd vccd _470_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[18\] _608_/Y mprj_logic_high_inst/HI[220] vssd vssd vccd
+ vccd la_oenb_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_9_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[75\]_A _537_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[93\]_B la_buf_enable\[93\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__570__A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_599_ la_oenb_mprj[9] vssd vssd vccd vccd _599_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y vssd vssd vccd vccd la_data_in_mprj[41]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[116\]_B user_to_mprj_in_gates\[116\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[84\]_B la_buf_enable\[84\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__480__A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__655__A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[75\]_B la_buf_enable\[75\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__390__A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[81\] la_iena_mprj[81] mprj_logic_high_inst/HI[411] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[81\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_522_ la_data_out_mprj[60] vssd vssd vccd vccd _522_/Y sky130_fd_sc_hd__inv_2
XANTENNA__565__A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_453_ mprj_dat_o_core[23] vssd vssd vccd vccd _453_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[45\] _507_/Y la_buf\[45\]/TE vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__einvp_8
X_384_ la_oenb_mprj[123] vssd vssd vccd vccd _384_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[117\] la_iena_mprj[117] mprj_logic_high_inst/HI[447] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[117\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[101\] _563_/Y la_buf\[101\]/TE vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_7_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y vssd vssd vccd vccd la_data_in_mprj[89]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] user_to_mprj_in_gates\[34\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[34\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__475__A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[57\]_B la_buf_enable\[57\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__385__A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[48\]_B la_buf_enable\[48\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[85\] _346_/Y mprj_logic_high_inst/HI[287] vssd vssd vccd
+ vccd la_oenb_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_2_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[108\] la_oenb_mprj[108] la_buf_enable\[108\]/B vssd vssd vccd vccd
+ la_buf\[108\]/TE sky130_fd_sc_hd__and2b_1
X_505_ la_data_out_mprj[43] vssd vssd vccd vccd _505_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[51\]_B mprj_logic_high_inst/HI[381] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[122\]_A_N la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_436_ mprj_dat_o_core[6] vssd vssd vccd vccd _436_/Y sky130_fd_sc_hd__inv_2
X_367_ la_oenb_mprj[106] vssd vssd vccd vccd _367_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[39\]_B la_buf_enable\[39\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[8\]_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[42\]_B mprj_logic_high_inst/HI[372] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[44\] la_iena_mprj[44] mprj_logic_high_inst/HI[374] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[44\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[33\]_B mprj_logic_high_inst/HI[363] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[22\] la_oenb_mprj[22] la_buf_enable\[22\]/B vssd vssd vccd vccd la_buf\[22\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[24\]_B mprj_logic_high_inst/HI[354] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_419_ mprj_adr_o_core[21] vssd vssd vccd vccd _419_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high_inst/HI[313] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[14\]_A _604_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] user_to_mprj_in_gates\[108\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[108\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[10\]_A _408_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[15\]_B mprj_logic_high_inst/HI[345] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high_inst/HI[212] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[118\] _379_/Y mprj_logic_high_inst/HI[320] vssd vssd vccd
+ vccd la_oenb_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_27_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[48\] _638_/Y mprj_logic_high_inst/HI[250] vssd vssd vccd
+ vccd la_oenb_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_1_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[2\]_B user_irq_ena_buf\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__573__A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_430 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[105] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y vssd vssd vccd vccd la_data_in_mprj[71]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__483__A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[33\]_TE mprj_logic_high_inst/HI[235] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[4\] _434_/Y mprj_dat_buf\[4\]/TE vssd vssd vccd vccd mprj_dat_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_316 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__393__A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_905 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__568__A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[80\]_A_N la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[23\]_A _453_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[75\] _537_/Y la_buf\[75\]/TE vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__einvp_8
XFILLER_1_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[95\]_A_N la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[33\]_A_N la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[48\]_A_N la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] user_to_mprj_in_gates\[64\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[64\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__478__A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__388__A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[79\]_TE mprj_logic_high_inst/HI[281] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_598_ la_oenb_mprj[8] vssd vssd vccd vccd _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y vssd vssd vccd vccd la_data_in_mprj[34]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[74\] la_iena_mprj[74] mprj_logic_high_inst/HI[404] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[74\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[100\] _361_/Y mprj_logic_high_inst/HI[302] vssd vssd vccd
+ vccd la_oenb_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_6_2291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[30\] _620_/Y mprj_logic_high_inst/HI[232] vssd vssd vccd
+ vccd la_oenb_core[30] sky130_fd_sc_hd__einvp_8
XFILLER_18_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_521_ la_data_out_mprj[59] vssd vssd vccd vccd _521_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[52\] la_oenb_mprj[52] la_buf_enable\[52\]/B vssd vssd vccd vccd la_buf\[52\]/TE
+ sky130_fd_sc_hd__and2b_1
X_452_ mprj_dat_o_core[22] vssd vssd vccd vccd _452_/Y sky130_fd_sc_hd__inv_2
X_383_ la_oenb_mprj[122] vssd vssd vccd vccd _383_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__581__A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[38\] _500_/Y la_buf\[38\]/TE vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_29_2248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2088 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] user_to_mprj_in_gates\[27\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[27\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__491__A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_A _406_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[78\] _339_/Y mprj_logic_high_inst/HI[280] vssd vssd vccd
+ vccd la_oenb_core[78] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[26\] _456_/Y mprj_dat_buf\[26\]/TE vssd vssd vccd vccd mprj_dat_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_24_2189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__576__A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_504_ la_data_out_mprj[42] vssd vssd vccd vccd _504_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_435_ mprj_dat_o_core[5] vssd vssd vccd vccd _435_/Y sky130_fd_sc_hd__inv_2
X_366_ la_oenb_mprj[105] vssd vssd vccd vccd _366_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[8\]_B mprj_logic_high_inst/HI[338] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[21\] _419_/Y mprj_adr_buf\[21\]/TE vssd vssd vccd vccd mprj_adr_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__486__A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[6\] la_oenb_mprj[6] la_buf_enable\[6\]/B vssd vssd vccd vccd la_buf\[6\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__396__A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_406 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[37\] la_iena_mprj[37] mprj_logic_high_inst/HI[367] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[37\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[15\] la_oenb_mprj[15] la_buf_enable\[15\]/B vssd vssd vccd vccd la_buf\[15\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[120\] la_oenb_mprj[120] la_buf_enable\[120\]/B vssd vssd vccd vccd
+ la_buf\[120\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_418_ mprj_adr_o_core[20] vssd vssd vccd vccd _418_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_349_ la_oenb_mprj[88] vssd vssd vccd vccd _349_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] user_to_mprj_in_gates\[94\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[94\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[121\]_A_N la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_2277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[20\] _482_/Y la_buf\[20\]/TE vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__einvp_8
XFILLER_8_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y vssd vssd vccd vccd la_data_in_mprj[64]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] user_to_mprj_in_gates\[120\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[120\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[110\]_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[60\] _650_/Y mprj_logic_high_inst/HI[262] vssd vssd vccd
+ vccd la_oenb_core[60] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[82\] la_oenb_mprj[82] la_buf_enable\[82\]/B vssd vssd vccd vccd la_buf\[82\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high_inst/HI[303] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__584__A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[68\] _530_/Y la_buf\[68\]/TE vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__einvp_8
XFILLER_16_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[101\]_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[124\] _586_/Y la_buf\[124\]/TE vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_6_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] user_to_mprj_in_gates\[57\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[57\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__494__A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_1_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1814 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high_inst/HI[326] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[90\]_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__579__A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[81\]_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_597_ la_oenb_mprj[7] vssd vssd vccd vccd _597_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y vssd vssd vccd vccd la_data_in_mprj[27]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__489__A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[72\]_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[8\]_B la_buf_enable\[8\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[94\]_A_N la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high_inst/HI[248] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__399__A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[67\] la_iena_mprj[67] mprj_logic_high_inst/HI[397] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[67\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_520_ la_data_out_mprj[58] vssd vssd vccd vccd _520_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[63\]_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[5\] _595_/Y mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd la_oenb_core[5] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[23\] _613_/Y mprj_logic_high_inst/HI[225] vssd vssd vccd
+ vccd la_oenb_core[23] sky130_fd_sc_hd__einvp_8
X_451_ mprj_dat_o_core[21] vssd vssd vccd vccd _451_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[45\] la_oenb_mprj[45] la_buf_enable\[45\]/B vssd vssd vccd vccd la_buf\[45\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[32\]_A_N la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_382_ la_oenb_mprj[121] vssd vssd vccd vccd _382_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[47\]_A_N la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_2191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[10\]_TE mprj_dat_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[54\]_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_649_ la_oenb_mprj[59] vssd vssd vccd vccd _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[84\]_TE la_buf\[84\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[69\]_TE mprj_logic_high_inst/HI[271] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[45\]_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[19\] _449_/Y mprj_dat_buf\[19\]/TE vssd vssd vccd vccd mprj_dat_o_user[19]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[36\]_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_503_ la_data_out_mprj[41] vssd vssd vccd vccd _503_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_434_ mprj_dat_o_core[4] vssd vssd vccd vccd _434_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__592__A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[50\] _512_/Y la_buf\[50\]/TE vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__einvp_8
X_365_ la_oenb_mprj[104] vssd vssd vccd vccd _365_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[122\] la_iena_mprj[122] mprj_logic_high_inst/HI[452] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[122\]/B sky130_fd_sc_hd__and2_1
XFILLER_14_698 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_A _433_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[14\] _412_/Y mprj_adr_buf\[14\]/TE vssd vssd vccd vccd mprj_adr_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y vssd vssd vccd vccd la_data_in_mprj[94]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[27\]_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] user_to_mprj_in_gates\[1\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[1\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[18\]_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[90\] _351_/Y mprj_logic_high_inst/HI[292] vssd vssd vccd
+ vccd la_oenb_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_3_845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[83\]_A user_to_mprj_in_gates\[83\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[98\] _560_/Y la_buf\[98\]/TE vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[3\] la_iena_mprj[3] mprj_logic_high_inst/HI[333] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[3\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__587__A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[113\] la_oenb_mprj[113] la_buf_enable\[113\]/B vssd vssd vccd vccd
+ la_buf\[113\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_2048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_417_ mprj_adr_o_core[19] vssd vssd vccd vccd _417_/Y sky130_fd_sc_hd__inv_2
X_348_ la_oenb_mprj[87] vssd vssd vccd vccd _348_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[110\]_A _572_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] user_to_mprj_in_gates\[87\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[87\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__497__A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[101\]_A _563_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y vssd vssd vccd vccd la_data_in_mprj[1]
+ sky130_fd_sc_hd__inv_8
XFILLER_31_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_281 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_454 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[13\] _475_/Y la_buf\[13\]/TE vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__einvp_8
Xla_buf\[9\] _471_/Y la_buf\[9\]/TE vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_3_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[6\] _404_/Y mprj_adr_buf\[6\]/TE vssd vssd vccd vccd mprj_adr_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_21_1982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y vssd vssd vccd vccd la_data_in_mprj[57]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_981 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[20\]_A _482_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] user_to_mprj_in_gates\[113\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[113\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_22_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[87\]_A _549_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[110\]_B mprj_logic_high_inst/HI[440] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[97\] la_iena_mprj[97] mprj_logic_high_inst/HI[427] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[97\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[123\] _384_/Y mprj_logic_high_inst/HI[325] vssd vssd vccd
+ vccd la_oenb_core[123] sky130_fd_sc_hd__einvp_8
XFILLER_5_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[53\] _643_/Y mprj_logic_high_inst/HI[255] vssd vssd vccd
+ vccd la_oenb_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_5_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[75\] la_oenb_mprj[75] la_buf_enable\[75\]/B vssd vssd vccd vccd la_buf\[75\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[101\]_B mprj_logic_high_inst/HI[431] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[96\]_B la_buf_enable\[96\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[117\] _579_/Y la_buf\[117\]/TE vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[110] sky130_fd_sc_hd__inv_8
XANTENNA_la_buf_enable\[20\]_B la_buf_enable\[20\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_B user_to_mprj_in_gates\[119\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[69\]_A _531_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_888 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[87\]_B la_buf_enable\[87\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[120\]_A_N la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[11\]_B la_buf_enable\[11\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2266 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[9\]_TE la_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[90\]_B mprj_logic_high_inst/HI[420] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_25_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[12\] la_iena_mprj[12] mprj_logic_high_inst/HI[342] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[12\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[78\]_B la_buf_enable\[78\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[80\] _542_/Y la_buf\[80\]/TE vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__einvp_8
XFILLER_29_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__595__A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_596_ la_oenb_mprj[6] vssd vssd vccd vccd _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[69\]_B la_buf_enable\[69\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_582 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[72\]_B mprj_logic_high_inst/HI[402] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_26_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_2063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[63\]_B mprj_logic_high_inst/HI[393] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_450_ mprj_dat_o_core[20] vssd vssd vccd vccd _450_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_313 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[16\] _606_/Y mprj_logic_high_inst/HI[218] vssd vssd vccd
+ vccd la_oenb_core[16] sky130_fd_sc_hd__einvp_8
X_381_ la_oenb_mprj[120] vssd vssd vccd vccd _381_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[38\] la_oenb_mprj[38] la_buf_enable\[38\]/B vssd vssd vccd vccd la_buf\[38\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[54\]_B mprj_logic_high_inst/HI[384] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_17_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_648_ la_oenb_mprj[58] vssd vssd vccd vccd _648_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_579_ la_data_out_mprj[117] vssd vssd vccd vccd _579_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[114\]_TE mprj_logic_high_inst/HI[316] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_917 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[45\]_B mprj_logic_high_inst/HI[375] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high_inst/HI[215] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_A _429_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[36\]_B mprj_logic_high_inst/HI[366] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_502_ la_data_out_mprj[40] vssd vssd vccd vccd _502_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_433_ mprj_dat_o_core[3] vssd vssd vccd vccd _433_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[43\] _505_/Y la_buf\[43\]/TE vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__einvp_8
X_364_ la_oenb_mprj[103] vssd vssd vccd vccd _364_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[115\] la_iena_mprj[115] mprj_logic_high_inst/HI[445] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[115\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1851 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y vssd vssd vccd vccd la_data_in_mprj[87]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_adr_buf\[22\]_A _420_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[27\]_B mprj_logic_high_inst/HI[357] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] user_to_mprj_in_gates\[32\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[32\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high_inst/HI[238] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[93\]_A_N la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[31\]_A_N la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[46\]_A_N la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[18\]_B mprj_logic_high_inst/HI[348] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[83\] _344_/Y mprj_logic_high_inst/HI[285] vssd vssd vccd
+ vccd la_oenb_core[83] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[31\] _461_/Y mprj_dat_buf\[31\]/TE vssd vssd vccd vccd mprj_dat_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[106\] la_oenb_mprj[106] la_buf_enable\[106\]/B vssd vssd vccd vccd
+ la_buf\[106\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_18_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1615 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_416_ mprj_adr_o_core[18] vssd vssd vccd vccd _416_/Y sky130_fd_sc_hd__inv_2
X_347_ la_oenb_mprj[86] vssd vssd vccd vccd _347_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_183 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[42\] la_iena_mprj[42] mprj_logic_high_inst/HI[372] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[42\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[20\] la_oenb_mprj[20] la_buf_enable\[20\]/B vssd vssd vccd vccd la_buf\[20\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__598__A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[26\]_A _456_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[17\]_A _447_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] user_to_mprj_in_gates\[106\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[106\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[116\] _377_/Y mprj_logic_high_inst/HI[318] vssd vssd vccd
+ vccd la_oenb_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_0_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[46\] _636_/Y mprj_logic_high_inst/HI[248] vssd vssd vccd
+ vccd la_oenb_core[46] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[68\] la_oenb_mprj[68] la_buf_enable\[68\]/B vssd vssd vccd vccd la_buf\[68\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_18_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[14\]_TE mprj_adr_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[103] sky130_fd_sc_hd__inv_8
XFILLER_19_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_dat_buf\[2\] _432_/Y mprj_dat_buf\[2\]/TE vssd vssd vccd vccd mprj_dat_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[110\]_B la_buf_enable\[110\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[73\] _535_/Y la_buf\[73\]/TE vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__einvp_8
XFILLER_38_2263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[101\]_B la_buf_enable\[101\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_595_ la_oenb_mprj[5] vssd vssd vccd vccd _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_594 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] user_to_mprj_in_gates\[62\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[62\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high_inst/HI[294] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_380_ la_oenb_mprj[119] vssd vssd vccd vccd _380_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_647_ la_oenb_mprj[57] vssd vssd vccd vccd _647_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_578_ la_data_out_mprj[116] vssd vssd vccd vccd _578_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y vssd vssd vccd vccd la_data_in_mprj[32]
+ sky130_fd_sc_hd__inv_8
XFILLER_31_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
.ends

