magic
tech sky130A
magscale 1 2
timestamp 1665590664
<< metal1 >>
rect 536 4 578 96
rect 606 4 648 96
rect 678 7 714 100
rect 742 7 788 100
<< metal2 >>
rect 20 -168 48 138
<< metal3 >>
rect -666 -1088 -2 -430
rect 78 -668 150 -508
<< metal4 >>
rect 516 -573 738 -440
rect 566 -652 738 -573
rect 821 -621 1219 -184
rect 516 -814 738 -652
<< rm5 >>
rect 821 -621 1219 -184
<< labels >>
flabel space -22 -322 -22 -322 0 FreeSans 320 0 0 0 Wide_spacing_rule
flabel space 612 -322 612 -322 0 FreeSans 320 0 0 0 Notch_rule
flabel space 614 228 614 228 0 FreeSans 320 0 0 0 Spacing_rule
flabel space 48 230 48 230 0 FreeSans 320 0 0 0 Width_rule
flabel space 604 -240 604 -240 0 FreeSans 320 0 0 0 Exercise_1d
flabel space 16 -244 16 -244 0 FreeSans 320 0 0 0 Exercise_1c
flabel space 608 296 608 296 0 FreeSans 320 0 0 0 Exercise_1b
flabel space 24 304 24 304 0 FreeSans 320 0 0 0 Exercise_1a
<< end >>
