magic
tech sky130A
timestamp 1665578704
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1665578704
transform 1 0 220 0 1 -1
box -19 -24 65 296
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1665578704
transform 1 0 -10 0 1 -1
box -19 -24 249 296
<< end >>
