* NGSPICE file created from inverter.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_BZBQCZ a_n173_n150# a_n78_n150# a_63_n238# a_n129_n238#
+ w_n311_n360# a_114_n150# a_18_n150# a_n33_172#
X0 a_114_n150# a_63_n238# a_18_n150# w_n311_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=180000u
X1 a_n78_n150# a_n129_n238# a_n173_n150# w_n311_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=180000u
X2 a_18_n150# a_n33_172# a_n78_n150# w_n311_n360# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=180000u
.ends

.subckt sky130_fd_pr__pfet_01v8_UTJYZV VSUBS a_n33_131# w_n311_n319# a_114_n100# a_63_n197#
+ a_18_n100# a_n129_n197# a_n173_n100# a_n78_n100#
X0 a_18_n100# a_n33_131# a_n78_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X1 a_114_n100# a_63_n197# a_18_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
X2 a_n78_n100# a_n129_n197# a_n173_n100# w_n311_n319# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=180000u
.ends

.subckt inverter in out vdd vss
XXM1 out vss in in vss vss out in sky130_fd_pr__nfet_01v8_BZBQCZ
XXM2 vss in vdd vdd in out in out vdd sky130_fd_pr__pfet_01v8_UTJYZV
.ends

